  
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[8]string"   p  0go.weak.type.**[8]string   �  type.[8]string   �8go.string.hdr."*[8]ast.Node"                       0go.string."*[8]ast.Node"   �0go.string."*[8]ast.Node"    *[8]ast.Node  � type.*[8]"".Node �  �              t.�a 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."*[8]ast.Node"   p  2go.weak.type.**[8]"".Node   �  type.[8]"".Node   �@go.string.hdr."*[8]interface {}"                       8go.string."*[8]interface {}"   �8go.string."*[8]interface {}" 0  "*[8]interface {}  �*type.*[8]interface {} �  �              �aK 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[8]interface {}"   p  <go.weak.type.**[8]interface {}   �  (type.[8]interface {}   �4go.string.hdr."*[7]string"             
          ,go.string."*[7]string"   �,go.string."*[7]string"    *[7]string  �type.*[7]string �  �              �Ϳ 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[7]string"   p  0go.weak.type.**[7]string   �  type.[7]string   �0go.string.hdr."go/token"                       (go.string."go/token"   �(go.string."go/token"    go/token  �.go.importpath.go/token.                       (go.string."go/token"   �&go.string.hdr."fmt"                       go.string."fmt"   �go.string."fmt"   fmt  �$go.importpath.fmt.                       go.string."fmt"   �.go.string.hdr."strconv"                       &go.string."strconv"   �&go.string."strconv"   strconv  �,go.importpath.strconv.                       &go.string."strconv"   �(go.string.hdr."sort"                        go.string."sort"   � go.string."sort"   
sort  �&go.importpath.sort.                        go.string."sort"   �.go.string.hdr."strings"                       &go.string."strings"   �&go.string."strings"   strings  �,go.importpath.strings.                       &go.string."strings"   �$go.string.hdr."io"                       go.string."io"   �go.string."io"   io  �"go.importpath.io.                       go.string."io"   �8go.string.hdr."unicode/utf8"                       0go.string."unicode/utf8"   �0go.string."unicode/utf8"    unicode/utf8  �6go.importpath.unicode/utf8.                       0go.string."unicode/utf8"   �.go.string.hdr."unicode"                       &go.string."unicode"   �&go.string."unicode"   unicode  �,go.importpath.unicode.                       &go.string."unicode"   �*go.string.hdr."bytes"                       "go.string."bytes"   �"go.string."bytes"   bytes  �(go.importpath.bytes.                       "go.string."bytes"   �$go.string.hdr."os"                       go.string."os"   �go.string."os"   os  �"go.importpath.os.                       go.string."os"   �.go.string.hdr."reflect"                       &go.string."reflect"   �&go.string."reflect"   reflect  �,go.importpath.reflect.                       &go.string."reflect"   �4go.string.hdr."go/scanner"             
          ,go.string."go/scanner"   �,go.string."go/scanner"    go/scanner  �2go.importpath.go/scanner.             
          ,go.string."go/scanner"   �0type..hash."".Comment·f              *type..hash."".Comment   �,type..eq."".Comment·f              &type..eq."".Comment   �0type..hash.[10]string·f              *type..hash.[10]string   �,type..eq.[10]string·f              &type..eq.[10]string   �."".(*ObjKind).String·f              ("".(*ObjKind).String   �.type..hash."".Object·f              (type..hash."".Object   �*type..eq."".Object·f              $type..eq."".Object   �,type..hash."".Ident·f              &type..hash."".Ident   �(type..eq."".Ident·f              "type..eq."".Ident   �"".Expr.End·f              "".Expr.End   �"".Expr.Pos·f              "".Expr.Pos   �&"".Expr.exprNode·f               "".Expr.exprNode   �2type..hash."".BasicLit·f              ,type..hash."".BasicLit   �.type..eq."".BasicLit·f              (type..eq."".BasicLit   �2type..hash."".Ellipsis·f              ,type..hash."".Ellipsis   �.type..eq."".Ellipsis·f              (type..eq."".Ellipsis   �"".Stmt.End·f              "".Stmt.End   �"".Stmt.Pos·f              "".Stmt.Pos   �&"".Stmt.stmtNode·f               "".Stmt.stmtNode   �4type..hash."".ParenExpr·f              .type..hash."".ParenExpr   �0type..eq."".ParenExpr·f              *type..eq."".ParenExpr   �:type..hash."".SelectorExpr·f              4type..hash."".SelectorExpr   �6type..eq."".SelectorExpr·f              0type..eq."".SelectorExpr   �4type..hash."".IndexExpr·f              .type..hash."".IndexExpr   �0type..eq."".IndexExpr·f              *type..eq."".IndexExpr   �4type..hash."".SliceExpr·f              .type..hash."".SliceExpr   �0type..eq."".SliceExpr·f              *type..eq."".SliceExpr   �>type..hash."".TypeAssertExpr·f              8type..hash."".TypeAssertExpr   �:type..eq."".TypeAssertExpr·f              4type..eq."".TypeAssertExpr   �2type..hash."".StarExpr·f              ,type..hash."".StarExpr   �.type..eq."".StarExpr·f              (type..eq."".StarExpr   �4type..hash."".UnaryExpr·f              .type..hash."".UnaryExpr   �0type..eq."".UnaryExpr·f              *type..eq."".UnaryExpr   �6type..hash."".BinaryExpr·f              0type..hash."".BinaryExpr   �2type..eq."".BinaryExpr·f              ,type..eq."".BinaryExpr   �:type..hash."".KeyValueExpr·f              4type..hash."".KeyValueExpr   �6type..eq."".KeyValueExpr·f              0type..eq."".KeyValueExpr   �4type..hash."".ArrayType·f              .type..hash."".ArrayType   �0type..eq."".ArrayType·f              *type..eq."".ArrayType   �6type..hash."".StructType·f              0type..hash."".StructType   �2type..eq."".StructType·f              ,type..eq."".StructType   �<type..hash."".InterfaceType·f              6type..hash."".InterfaceType   �8type..eq."".InterfaceType·f              2type..eq."".InterfaceType   �0type..hash."".MapType·f              *type..hash."".MapType   �,type..eq."".MapType·f              &type..eq."".MapType   �2type..hash."".ChanType·f              ,type..hash."".ChanType   �.type..eq."".ChanType·f              (type..eq."".ChanType   �"".Decl.End·f              "".Decl.End   �"".Decl.Pos·f              "".Decl.Pos   �&"".Decl.declNode·f               "".Decl.declNode   �4type..hash."".EmptyStmt·f              .type..hash."".EmptyStmt   �0type..eq."".EmptyStmt·f              *type..eq."".EmptyStmt   �8type..hash."".LabeledStmt·f              2type..hash."".LabeledStmt   �4type..eq."".LabeledStmt·f              .type..eq."".LabeledStmt   �2type..hash."".SendStmt·f              ,type..hash."".SendStmt   �.type..eq."".SendStmt·f              (type..eq."".SendStmt   �6type..hash."".IncDecStmt·f              0type..hash."".IncDecStmt   �2type..eq."".IncDecStmt·f              ,type..eq."".IncDecStmt   �.type..hash."".IfStmt·f              (type..hash."".IfStmt   �*type..eq."".IfStmt·f              $type..eq."".IfStmt   �6type..hash."".SwitchStmt·f              0type..hash."".SwitchStmt   �2type..eq."".SwitchStmt·f              ,type..eq."".SwitchStmt   �>type..hash."".TypeSwitchStmt·f              8type..hash."".TypeSwitchStmt   �:type..eq."".TypeSwitchStmt·f              4type..eq."".TypeSwitchStmt   �0type..hash."".ForStmt·f              *type..hash."".ForStmt   �,type..eq."".ForStmt·f              &type..eq."".ForStmt   �4type..hash."".RangeStmt·f              .type..hash."".RangeStmt   �0type..eq."".RangeStmt·f              *type..eq."".RangeStmt   �2type..hash."".TypeSpec·f              ,type..hash."".TypeSpec   �.type..eq."".TypeSpec·f              (type..eq."".TypeSpec   �"".Spec.End·f              "".Spec.End   �"".Spec.Pos·f              "".Spec.Pos   �&"".Spec.specNode·f               "".Spec.specNode   �.type..hash.[8]string·f              (type..hash.[8]string   �*type..eq.[8]string·f              $type..eq.[8]string   �$"".(*byPos).Len·f              "".(*byPos).Len   �&"".(*byPos).Less·f               "".(*byPos).Less   �&"".(*byPos).Swap·f               "".(*byPos).Swap   �"".Node.End·f              "".Node.End   �"".Node.Pos·f              "".Node.Pos   �0type..hash.[8]"".Node·f              *type..hash.[8]"".Node   �,type..eq.[8]"".Node·f              &type..eq.[8]"".Node   �<"".(*CommentMap).addComment·f              6"".(*CommentMap).addComment   �4"".(*CommentMap).Update·f              ."".(*CommentMap).Update   �4"".(*CommentMap).Filter·f              ."".(*CommentMap).Filter   �8"".(*CommentMap).Comments·f              2"".(*CommentMap).Comments   �4"".(*CommentMap).String·f              ."".(*CommentMap).String   �."".(*byInterval).Len·f              ("".(*byInterval).Len   �0"".(*byInterval).Less·f              *"".(*byInterval).Less   �0"".(*byInterval).Swap·f              *"".(*byInterval).Swap   �:type..hash.[1]interface {}·f              4type..hash.[1]interface {}   �6type..eq.[1]interface {}·f              0type..eq.[1]interface {}   �:type..hash.[3]interface {}·f              4type..hash.[3]interface {}   �6type..eq.[3]interface {}·f              0type..eq.[3]interface {}   �2"".(*byImportSpec).Len·f              ,"".(*byImportSpec).Len   �4"".(*byImportSpec).Swap·f              ."".(*byImportSpec).Swap   �4"".(*byImportSpec).Less·f              ."".(*byImportSpec).Less   �2"".(*byCommentPos).Len·f              ,"".(*byCommentPos).Len   �4"".(*byCommentPos).Swap·f              ."".(*byCommentPos).Swap   �4"".(*byCommentPos).Less·f              ."".(*byCommentPos).Less   �:type..hash.[8]interface {}·f              4type..hash.[8]interface {}   �6type..eq.[8]interface {}·f              0type..eq.[8]interface {}   �:type..hash.[2]interface {}·f              4type..hash.[2]interface {}   �6type..eq.[2]interface {}·f              0type..eq.[2]interface {}   �&"".Visitor.Visit·f               "".Visitor.Visit   �0"".(*inspector).Visit·f              *"".(*inspector).Visit   �.type..hash.[7]string·f              (type..hash.[7]string   �*type..eq.[7]string·f              $type..eq.[7]string   ��go13ld       usr/local/go/pkg/linux_amd64/go/build.a                                                             0100644 0000000 0000000 00001327632 13101127332 016345  0                                                                                                    ustar 00                                                                0000000 0000000                                                                                                                                                                        !<arch>
__.PKGDEF       0           0     0     644     16693     `
go object linux amd64 go1.6.4 X:none
build id "23f3739002c9f2b861ac9117ef7aa0e5f75cb85f"

$$
package build
	import runtime "runtime"
	import bytes "bytes"
	import errors "errors"
	import io "io"
	import utf8 "unicode/utf8"
	import unicode "unicode"
	import fmt "fmt"
	import strconv "strconv"
	import os "os"
	import ast "go/ast"
	import token "go/token"
	import sort "sort"
	import strings "strings"
	import doc "go/doc"
	import path "path"
	import parser "go/parser"
	import ioutil "io/ioutil"
	import filepath "path/filepath"
	import log "log"
	import bufio "bufio"
	import time "time" // indirect
	type @"time".zone struct { @"time".name string; @"time".offset int; @"time".isDST bool }
	type @"time".zoneTrans struct { @"time".when int64; @"time".index uint8; @"time".isstd bool; @"time".isutc bool }
	type @"time".Location struct { @"time".name string; @"time".zone []@"time".zone; @"time".tx []@"time".zoneTrans; @"time".cacheStart int64; @"time".cacheEnd int64; @"time".cacheZone *@"time".zone }
	func (@"time".l·2 *@"time".Location "esc:0x22") String () (? string)
	func (@"time".l·2 *@"time".Location "esc:0x1") @"time".firstZoneUsed () (? bool)
	func (@"time".l·2 *@"time".Location "esc:0x12") @"time".get () (? *@"time".Location)
	func (@"time".l·6 *@"time".Location "esc:0x32") @"time".lookup (@"time".sec·7 int64) (@"time".name·1 string, @"time".offset·2 int, @"time".isDST·3 bool, @"time".start·4 int64, @"time".end·5 int64)
	func (@"time".l·2 *@"time".Location "esc:0x1") @"time".lookupFirstZone () (? int)
	func (@"time".l·4 *@"time".Location "esc:0x1") @"time".lookupName (@"time".name·5 string "esc:0x1", @"time".unix·6 int64) (@"time".offset·1 int, @"time".isDST·2 bool, @"time".ok·3 bool)
	type @"time".Duration int64
	func (@"time".d·2 @"time".Duration) Hours () (? float64) { var @"time".hour·3 @"time".Duration; ; @"time".hour·3 = @"time".d·2 / @"time".Duration(0x34630b8a000); var @"time".nsec·4 @"time".Duration; ; @"time".nsec·4 = @"time".d·2 % @"time".Duration(0x34630b8a000); return float64(@"time".hour·3) + float64(@"time".nsec·4) * float64(8190022623310637111963488201822504381538623676021880892417778544696899264837610290203272971060556344039023584360473938041055625214280336402169897364226048p-553) }
	func (@"time".d·2 @"time".Duration) Minutes () (? float64) { var @"time".min·3 @"time".Duration; ; @"time".min·3 = @"time".d·2 / @"time".Duration(0xdf8475800); var @"time".nsec·4 @"time".Duration; ; @"time".nsec·4 = @"time".d·2 % @"time".Duration(0xdf8475800); return float64(@"time".min·3) + float64(@"time".nsec·4) * float64(7678146209353722106395056769533233877065564876941352542109479049699919628723768656821910653339403201031675627614471533358284117434246264392176261853609984p-547) }
	func (@"time".d·2 @"time".Duration) Nanoseconds () (? int64) { return int64(@"time".d·2) }
	func (@"time".d·2 @"time".Duration) Seconds () (? float64) { var @"time".sec·3 @"time".Duration; ; @"time".sec·3 = @"time".d·2 / @"time".Duration(0x3b9aca00); var @"time".nsec·4 @"time".Duration; ; @"time".nsec·4 = @"time".d·2 % @"time".Duration(0x3b9aca00); return float64(@"time".sec·3) + float64(@"time".nsec·4) * float64(7198262071269114660816079141112770740375861891461678802759824945047098083990024106014198994535558872472104883612039846078596891298747423852523262413111296p-541) }
	func (@"time".d·2 @"time".Duration) String () (? string)
	type @"time".Month int
	func (@"time".m·2 @"time".Month) String () (? string) { return @"time".months[@"time".m·2 - @"time".Month(0x1)] }
	type @"time".Weekday int
	func (@"time".d·2 @"time".Weekday) String () (? string) { return @"time".days[@"time".d·2] }
	type @"time".Time struct { @"time".sec int64; @"time".nsec int32; @"time".loc *@"time".Location }
	func (@"time".t·2 @"time".Time "esc:0x12") Add (@"time".d·3 @"time".Duration) (? @"time".Time) { @"time".t·2.@"time".sec += int64(@"time".d·3 / @"time".Duration(0x3b9aca00)); var @"time".nsec·4 int32; ; @"time".nsec·4 = int32(@"time".t·2.@"time".nsec) + int32(@"time".d·3 % @"time".Duration(0x3b9aca00)); if @"time".nsec·4 >= int32(0x3b9aca00) { @"time".t·2.@"time".sec++; @"time".nsec·4 -= int32(0x3b9aca00) } else { if @"time".nsec·4 < int32(0x0) { @"time".t·2.@"time".sec--; @"time".nsec·4 += int32(0x3b9aca00) } }; @"time".t·2.@"time".nsec = @"time".nsec·4; return @"time".t·2 }
	func (@"time".t·2 @"time".Time "esc:0x12") AddDate (@"time".years·3 int, @"time".months·4 int, @"time".days·5 int) (? @"time".Time)
	func (@"time".t·2 @"time".Time "esc:0x1") After (@"time".u·3 @"time".Time "esc:0x1") (? bool) { return @"time".t·2.@"time".sec > @"time".u·3.@"time".sec || @"time".t·2.@"time".sec == @"time".u·3.@"time".sec && @"time".t·2.@"time".nsec > @"time".u·3.@"time".nsec }
	func (@"time".t·2 @"time".Time "esc:0x9") AppendFormat (@"time".b·3 []byte "esc:0x1a", @"time".layout·4 string "esc:0x9") (? []byte)
	func (@"time".t·2 @"time".Time "esc:0x1") Before (@"time".u·3 @"time".Time "esc:0x1") (? bool) { return @"time".t·2.@"time".sec < @"time".u·3.@"time".sec || @"time".t·2.@"time".sec == @"time".u·3.@"time".sec && @"time".t·2.@"time".nsec < @"time".u·3.@"time".nsec }
	func (@"time".t·4 @"time".Time "esc:0x1") Clock () (@"time".hour·1 int, @"time".min·2 int, @"time".sec·3 int)
	func (@"time".t·4 @"time".Time "esc:0x1") Date () (@"time".year·1 int, @"time".month·2 @"time".Month, @"time".day·3 int)
	func (@"time".t·2 @"time".Time "esc:0x1") Day () (? int)
	func (@"time".t·2 @"time".Time "esc:0x1") Equal (@"time".u·3 @"time".Time "esc:0x1") (? bool) { return @"time".t·2.@"time".sec == @"time".u·3.@"time".sec && @"time".t·2.@"time".nsec == @"time".u·3.@"time".nsec }
	func (@"time".t·2 @"time".Time "esc:0x9") Format (@"time".layout·3 string "esc:0x9") (? string)
	func (@"time".t·2 *@"time".Time "esc:0x1") GobDecode (@"time".data·3 []byte "esc:0x1") (? error)
	func (@"time".t·3 @"time".Time "esc:0x1") GobEncode () (? []byte, ? error)
	func (@"time".t·2 @"time".Time "esc:0x1") Hour () (? int)
	func (@"time".t·3 @"time".Time "esc:0x1") ISOWeek () (@"time".year·1 int, @"time".week·2 int)
	func (@"time".t·2 @"time".Time "esc:0x12") In (@"time".loc·3 *@"time".Location "esc:0x12") (? @"time".Time)
	func (@"time".t·2 @"time".Time "esc:0x1") IsZero () (? bool) { return @"time".t·2.@"time".sec == int64(0x0) && @"time".t·2.@"time".nsec == int32(0x0) }
	func (@"time".t·2 @"time".Time "esc:0x12") Local () (? @"time".Time) { @"time".t·2.@"time".loc = @"time".Local; return @"time".t·2 }
	func (@"time".t·2 @"time".Time "esc:0x12") Location () (? *@"time".Location) { var @"time".l·3 *@"time".Location; ; @"time".l·3 = @"time".t·2.@"time".loc; if @"time".l·3 == nil { @"time".l·3 = @"time".UTC }; return @"time".l·3 }
	func (@"time".t·3 @"time".Time "esc:0x1") MarshalBinary () (? []byte, ? error)
	func (@"time".t·3 @"time".Time "esc:0x9") MarshalJSON () (? []byte, ? error)
	func (@"time".t·3 @"time".Time "esc:0x9") MarshalText () (? []byte, ? error)
	func (@"time".t·2 @"time".Time "esc:0x1") Minute () (? int)
	func (@"time".t·2 @"time".Time "esc:0x1") Month () (? @"time".Month)
	func (@"time".t·2 @"time".Time "esc:0x1") Nanosecond () (? int) { return int(@"time".t·2.@"time".nsec) }
	func (@"time".t·2 @"time".Time "esc:0x12") Round (@"time".d·3 @"time".Duration) (? @"time".Time)
	func (@"time".t·2 @"time".Time "esc:0x1") Second () (? int)
	func (@"time".t·2 @"time".Time "esc:0x9") String () (? string)
	func (@"time".t·2 @"time".Time "esc:0x1") Sub (@"time".u·3 @"time".Time "esc:0x1") (? @"time".Duration)
	func (@"time".t·2 @"time".Time "esc:0x12") Truncate (@"time".d·3 @"time".Duration) (? @"time".Time)
	func (@"time".t·2 @"time".Time "esc:0x12") UTC () (? @"time".Time) { @"time".t·2.@"time".loc = @"time".UTC; return @"time".t·2 }
	func (@"time".t·2 @"time".Time "esc:0x1") Unix () (? int64) { return @"time".t·2.@"time".sec + int64(-0xe7791f700) }
	func (@"time".t·2 @"time".Time "esc:0x1") UnixNano () (? int64) { return (@"time".t·2.@"time".sec + int64(-0xe7791f700)) * int64(0x3b9aca00) + int64(@"time".t·2.@"time".nsec) }
	func (@"time".t·2 *@"time".Time "esc:0x1") UnmarshalBinary (@"time".data·3 []byte "esc:0x1") (? error)
	func (@"time".t·2 *@"time".Time "esc:0x1") UnmarshalJSON (@"time".data·3 []byte "esc:0x1") (@"time".err·1 error)
	func (@"time".t·2 *@"time".Time "esc:0x1") UnmarshalText (@"time".data·3 []byte "esc:0x1") (@"time".err·1 error)
	func (@"time".t·2 @"time".Time "esc:0x1") Weekday () (? @"time".Weekday)
	func (@"time".t·2 @"time".Time "esc:0x1") Year () (? int)
	func (@"time".t·2 @"time".Time "esc:0x1") YearDay () (? int)
	func (@"time".t·3 @"time".Time "esc:0x32") Zone () (@"time".name·1 string, @"time".offset·2 int)
	func (@"time".t·2 @"time".Time "esc:0x1") @"time".abs () (? uint64)
	func (@"time".t·5 @"time".Time "esc:0x1") @"time".date (@"time".full·6 bool) (@"time".year·1 int, @"time".month·2 @"time".Month, @"time".day·3 int, @"time".yday·4 int)
	func (@"time".t·4 @"time".Time "esc:0x32") @"time".locabs () (@"time".name·1 string, @"time".offset·2 int, @"time".abs·3 uint64)
	type @"os".FileMode uint32
	func (@"os".m·2 @"os".FileMode) IsDir () (? bool) { return @"os".m·2 & @"os".FileMode(0x80000000) != @"os".FileMode(0x0) }
	func (@"os".m·2 @"os".FileMode) IsRegular () (? bool) { return @"os".m·2 & @"os".FileMode(0x8f000000) == @"os".FileMode(0x0) }
	func (@"os".m·2 @"os".FileMode) Perm () (? @"os".FileMode) { return @"os".m·2 & @"os".FileMode(0x1ff) }
	func (@"os".m·2 @"os".FileMode) String () (? string)
	type @"os".FileInfo interface { IsDir() (? bool); ModTime() (? @"time".Time); Mode() (? @"os".FileMode); Name() (? string); Size() (? int64); Sys() (? interface {}) }
	type @"io".ReadCloser interface { Close() (? error); Read(@"io".p []byte) (@"io".n int, @"io".err error) }
	type @"go/token".Position struct { Filename string; Offset int; Line int; Column int }
	func (@"go/token".pos·2 *@"go/token".Position "esc:0x1") IsValid () (? bool) { return @"go/token".pos·2.Line > int(0x0) }
	func (@"go/token".pos·2 @"go/token".Position "esc:0x12") String () (? string)
	type @"".Package struct { Dir string; Name string; ImportComment string; Doc string; ImportPath string; Root string; SrcRoot string; PkgRoot string; PkgTargetRoot string; BinDir string; Goroot bool; PkgObj string; AllTags []string; ConflictDir string; GoFiles []string; CgoFiles []string; IgnoredGoFiles []string; InvalidGoFiles []string; CFiles []string; CXXFiles []string; MFiles []string; HFiles []string; SFiles []string; SwigFiles []string; SwigCXXFiles []string; SysoFiles []string; CgoCFLAGS []string; CgoCPPFLAGS []string; CgoCXXFLAGS []string; CgoLDFLAGS []string; CgoPkgConfig []string; Imports []string; ImportPos map[string][]@"go/token".Position; TestGoFiles []string; TestImports []string; TestImportPos map[string][]@"go/token".Position; XTestGoFiles []string; XTestImports []string; XTestImportPos map[string][]@"go/token".Position }
	func (@"".p·2 *@"".Package "esc:0x1") IsCommand () (? bool) { return @"".p·2.Name == string("main") }
	type @"".ImportMode uint
	type @"go/token".Pos int
	func (@"go/token".p·2 @"go/token".Pos) IsValid () (? bool) { return @"go/token".p·2 != @"go/token".Pos(0x0) }
	type @"go/ast".Comment struct { Slash @"go/token".Pos; Text string }
	func (@"go/ast".c·2 *@"go/ast".Comment "esc:0x1") End () (? @"go/token".Pos) { return @"go/token".Pos(int(@"go/ast".c·2.Slash) + len(@"go/ast".c·2.Text)) }
	func (@"go/ast".c·2 *@"go/ast".Comment "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".c·2.Slash }
	type @"go/ast".CommentGroup struct { List []*@"go/ast".Comment }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x1") End () (? @"go/token".Pos) { return @"go/ast".g·2.List[len(@"go/ast".g·2.List) - int(0x1)].End() }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".g·2.List[int(0x0)].Pos() }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x9") Text () (? string)
	type @"".Context struct { GOARCH string; GOOS string; GOROOT string; GOPATH string; CgoEnabled bool; UseAllFiles bool; Compiler string; BuildTags []string; ReleaseTags []string; InstallSuffix string; JoinPath func(@"".elem ...string) (? string); SplitPathList func(@"".list string) (? []string); IsAbsPath func(@"".path string) (? bool); IsDir func(@"".path string) (? bool); HasSubdir func(@"".root string, @"".dir string) (@"".rel string, @"".ok bool); ReadDir func(@"".dir string) (@"".fi []@"os".FileInfo, @"".err error); OpenFile func(@"".path string) (@"".r @"io".ReadCloser, @"".err error) }
	func (@"".ctxt·3 *@"".Context "esc:0x18a") Import (@"".path·4 string, @"".srcDir·5 string, @"".mode·6 @"".ImportMode) (? *@"".Package, ? error)
	func (@"".ctxt·3 *@"".Context "esc:0x18a") ImportDir (@"".dir·4 string, @"".mode·5 @"".ImportMode) (? *@"".Package, ? error)
	func (@"".ctxt·3 *@"".Context "esc:0x18a") MatchFile (@"".dir·4 string, @"".name·5 string) (@"".match·1 bool, @"".err·2 error)
	func (@"".ctxt·2 *@"".Context "esc:0x9") SrcDirs () (? []string)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".goodOSArchFile (@"".name·3 string, @"".allTags·4 map[string]bool "esc:0x1") (? bool)
	func (@"".ctxt·2 *@"".Context "esc:0x9") @"".gopath () (? []string)
	func (@"".ctxt·3 *@"".Context "esc:0x32") @"".hasSubdir (@"".root·4 string, @"".dir·5 string) (@"".rel·1 string, @"".ok·2 bool)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".isAbsPath (@"".path·3 string) (? bool)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".isDir (@"".path·3 string) (? bool)
	func (@"".ctxt·2 *@"".Context "esc:0x9") @"".isFile (@"".path·3 string) (? bool)
	func (@"".ctxt·2 *@"".Context "esc:0x32") @"".joinPath (@"".elem·3 ...string) (? string)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".match (@"".name·3 string, @"".allTags·4 map[string]bool "esc:0x1") (? bool)
	func (@"".ctxt·5 *@"".Context "esc:0x6c0a") @"".matchFile (@"".dir·6 string, @"".name·7 string, @"".returnImports·8 bool, @"".allTags·9 map[string]bool "esc:0x1") (@"".match·1 bool, @"".data·2 []byte, @"".filename·3 string, @"".err·4 error)
	func (@"".ctxt·3 *@"".Context "esc:0x1b2") @"".openFile (@"".path·4 string) (? @"io".ReadCloser, ? error)
	func (@"".ctxt·3 *@"".Context "esc:0x1b2") @"".readDir (@"".path·4 string) (? []@"os".FileInfo, ? error)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".saveCgo (@"".filename·3 string, @"".di·4 *@"".Package "esc:0x9", @"".cg·5 *@"go/ast".CommentGroup "esc:0x9") (? error)
	func (@"".ctxt·2 *@"".Context "esc:0x1") @"".shouldBuild (@"".content·3 []byte "esc:0x1", @"".allTags·4 map[string]bool "esc:0x1") (? bool)
	func (@"".ctxt·2 *@"".Context "esc:0x32") @"".splitPathList (@"".s·3 string) (? []string)
	var @"".Default @"".Context
	const @"".FindOnly @"".ImportMode = 0x1
	const @"".AllowBinary @"".ImportMode = 0x2
	const @"".ImportComment @"".ImportMode = 0x4
	const @"".IgnoreVendor @"".ImportMode = 0x8
	type @"".NoGoError struct { Dir string }
	func (@"".e·2 *@"".NoGoError "esc:0x1") Error () (? string) { return string("no buildable Go source files in ") + @"".e·2.Dir }
	type @"".MultiplePackageError struct { Dir string; Packages []string; Files []string }
	func (@"".e·2 *@"".MultiplePackageError "esc:0x9") Error () (? string)
	func @"".Import (@"".path·3 string, @"".srcDir·4 string, @"".mode·5 @"".ImportMode) (? *@"".Package, ? error)
	func @"".ImportDir (@"".dir·3 string, @"".mode·4 @"".ImportMode) (? *@"".Package, ? error)
	var @"".ToolDir string
	func @"".IsLocalImport (@"".path·2 string "esc:0x1") (? bool) { return @"".path·2 == string(".") || @"".path·2 == string("..") || @"strings".HasPrefix(@"".path·2, string("./")) || @"strings".HasPrefix(@"".path·2, string("../")) }
	func @"".ArchChar (@"".goarch·3 string "esc:0x1") (? string, ? error) { return string("?"), @"errors".New(string("architecture letter no longer used")) }
	func @"".init ()
	var @"time".months [12]string
	var @"time".days [7]string
	var @"time".Local *@"time".Location
	var @"time".UTC *@"time".Location
	func @"strings".HasPrefix (@"strings".s·2 string "esc:0x1", @"strings".prefix·3 string "esc:0x1") (? bool) { return len(@"strings".s·2) >= len(@"strings".prefix·3) && @"strings".s·2[int(0x0):len(@"strings".prefix·3)] == @"strings".prefix·3 }
	func @"errors".New (@"errors".text·2 string) (? error) { return (&@"errors".errorString{ @"errors".s:@"errors".text·2 }) }
	type @"errors".errorString struct { @"errors".s string }
	func (@"errors".e·2 *@"errors".errorString "esc:0x22") Error () (? string) { return @"errors".e·2.@"errors".s }

$$
 _go_.o          0           0     0     644     355811    `
go object linux amd64 go1.6.4 X:none

!
  go13ldbytes.aerrors.a
fmt.ago/ast.ago/doc.ago/parser.ago/token.aio.aio/ioutil.a
log.aos.apath.apath/filepath.aruntime.asort.astrconv.astrings.aunicode.aunicode/utf8.abufio.a �,"".(*Context).joinPath  �  �dH�%    H;a��   H��(H�t$8H�T$@H�L$H1�H�\$PH�\$XH�\$0H���   1�H9�t/H�4$H�T$H�L$H�H����H�L$H�D$ H�L$PH�D$XH��(�H�4$H�T$H�L$�    H�L$H�D$ H�L$PH�D$XH��(��    �V���������
      �       �  $path/filepath.Join   �  0runtime.morestack_noctxt   `P  "".autotmp_0001  type.string "".~r1 @type.string "".elem type.[]string "".ctxt   type.*"".Context P\OP+O � �2/, 
 YW Tgclocals·d98f60bd8519d0c68364b2a1d83af357 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�6"".(*Context).splitPathList  �  �dH�%    H;a��   H��(H�T$8H�L$@1�H�\$HH�\$PH�\$XH�\$0H���   1�H9�t4H�$H�L$H�H����H�T$H�L$H�D$ H�T$HH�L$PH�D$XH��(�H�$H�L$�    H�T$H�L$H�D$ H�T$HH�L$PH�D$XH��(��    �L���������������
      �       �  .path/filepath.SplitList   �  0runtime.morestack_noctxt   `P  "".autotmp_0003  type.[]string "".~r1 0type.[]string "".s type.string "".ctxt   type.*"".Context PaOP0O � �241 
 Tl Tgclocals·d98f60bd8519d0c68364b2a1d83af357 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�."".(*Context).isAbsPath  �  �dH�%    H;a��   H��hH�L$xH��$�   H�\$pH���   1�H9�t"H�$H�T$H�H�����\$��$�   H��h�H�L$HH�T$PH�=    H��   H9�|_H�T$0H9�wNH�L$(H9�u@H�L$XH�$H�D$`H�D$H�|$8H�|$H�D$@H�D$�    �\$ H�؈�$�   H��h�1����    1����    �����������������
      �       �  go.string."/"   �   runtime.eqstring   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0010  type.bool "".autotmp_0009  type.bool "".autotmp_0008 type.string "strings.prefix·3 _type.string strings.s·2 type.string *path/filepath.path·2 ?type.string "".~r1 0type.bool "".path type.string "".ctxt   type.*"".Context *�A��p��� � �$"�  F� Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·895d0569a38a56443b84805daa09d838   :$GOROOT/src/go/build/build.go�&"".(*Context).isDir  �  �dH�%    H;a��   H��PH�T$`H�L$hH�\$XH���   1�H9�tH�$H�L$H�H�����\$�\$pH��P�H�$H�L$�    H�T$H�L$H�D$ H�\$(H�\$HH�D$@H�� u"H�L$8H�$H�T$0H�Z ���\$�\$pH��P��D$p ���    �H�����������

      �       �  os.Stat   �       �  0runtime.morestack_noctxt   @�  "".autotmp_0012  type.bool "".err type.error 
"".fi ? type.os.FileInfo "".~r1 0type.bool "".path type.string "".ctxt   type.*"".Context *�;��S��� � �!'4	 
 C} Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�."".(*Context).hasSubdir  �	  �	dH�%    H;a�=  H��XH�|$hH�t$pH�T$xH��$�   1�1�H��$�   H��$�   H�\$`H���   1�H9�tFH�<$H�t$H�T$H�L$H�H����H�T$ H�L$(�\$0H��$�   H��$�   ��$�   H��X�H�<$H�t$H�T$H�L$�    H�\$ H��$�   H�\$(H��$�   �\$0�� ��$�   tH��X�H�\$hH�$H�\$pH�\$�    H�\$H�\$8H�\$H�\$@H�\$xH�$H��$�   H�\$�    H�\$H�\$HH�\$H�\$PH�\$8H�$H�\$@H�\$H�\$xH�\$H��$�   H�\$�    H�\$ H��$�   H�\$(H��$�   �\$0�� ��$�   tH��X�H�\$hH�$H�\$pH�\$H�\$HH�\$H�\$PH�\$�    H�\$ H��$�   H�\$(H��$�   �\$0�� ��$�   tH��X�H�\$8H�$H�\$@H�\$H�\$HH�\$H�\$PH�\$�    H�T$ H�L$(�\$0H��$�   H��$�   ��$�   H��X��    ����������
      �       �  "".hasSubdir   �  4path/filepath.EvalSymlinks   �  4path/filepath.EvalSymlinks   �  "".hasSubdir   �  "".hasSubdir   �  "".hasSubdir   �	  0runtime.morestack_noctxt   ��  "".autotmp_0016  type.bool "".autotmp_0015  type.string "".dirSym type.string "".rootSym ?type.string 
"".ok ptype.bool "".rel Ptype.string "".dir 0type.string "".root type.string "".ctxt   type.*"".Context F����G�����[��V� � 8�BFC,/ZWW+  n�C�@ Tgclocals·dd9ae044070cfdff36caf84fd74b60b9 Tgclocals·b4e92317a1ad7fa1f283390980fe4780   :$GOROOT/src/go/build/build.go�"".hasSubdir  �  �dH�%    H�D$�H;A��  H��   1�1�H��$�   H��$�   H��$�   H�$H��$�   H�\$�    L�T$L�L$L��$�   L�T$8L��$�   H�5    H�t$XH��   L�L$@H�D$`I9��(  L��H)�L��L9��  H)�M��H�� tM�H9���  L�D$xL�$H��$�   H�l$H�t$H�D$�    L��$�   L��$�   �\$ H��< uSH�$    L�T$xL�T$L��$�   L�L$H�    H�\$H�D$    �    H�\$(H��$�   H�\$0H��$�   H��$�   H�$H��$�   H�\$�    L�L$L�D$L��$�   L�L$HL��$�   H��$�   H�t$hH��$�   L�D$PH�D$pI9���   L9���   H9���   L�L$xL�$H��$�   H�D$H�t$H�D$�    L��$�   L��$�   �\$ H��< u"1�H��$�   H��$�   Ƅ$�    H�Ĉ   �H��$�   L��L9�wUH)�M��H�� tM�L�D$xL�$H��$�   H�l$�    H�D$H�L$H��$�   H��$�   Ƅ$�   H�Ĉ   ��    1��g����    1��Y���1��G����    1��9����    �1����
      �  &path/filepath.Clean   �  go.string."/"   �   runtime.eqstring   �  go.string."/"   �  *runtime.concatstring2   �  &path/filepath.Clean   �   runtime.eqstring   �	  *path/filepath.ToSlash   �
  $runtime.panicslice   �
  $runtime.panicslice   �
  $runtime.panicslice   �  0runtime.morestack_noctxt   p�  $"".autotmp_0032  type.bool "".autotmp_0030  type.string "".autotmp_0029  type.string "".autotmp_0028  type.int "".autotmp_0027  type.string "".autotmp_0026  type.int "".autotmp_0025  type.int "".autotmp_0024  type.int "".autotmp_0023  type.string "".autotmp_0022 type.string "strings.prefix·3 ?type.string strings.s·2 type.string "strings.suffix·3 _type.string strings.s·2 �type.string 
"".ok `type.bool "".rel @type.string "".dir  type.string "".root  type.string ,����d��1� � 4�3(�S(�"l  L� Tgclocals·12ab5efd4c34ee1072eaafe77351d565 Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c   :$GOROOT/src/go/build/build.go�*"".(*Context).readDir  �  �dH�%    H;a��   H��8H�T$HH�L$P1�H�\$XH�\$`H�\$h1�H�\$pH�\$xH�\$@H���   1�H9�tHH�$H�L$H�H����H�t$H�l$H�T$ H�L$(H�D$0H�t$XH�l$`H�T$hH�L$pH�D$xH��8�H�$H�L$�    H�t$H�l$H�T$ H�L$(H�D$0H�t$XH�l$`H�T$hH�L$pH�D$xH��8��    ������������
      �       �  "io/ioutil.ReadDir   �  0runtime.morestack_noctxt   �p  "".autotmp_0036  type.error "".autotmp_0035  $type.[]os.FileInfo "".~r2 `type.error "".~r1 0$type.[]os.FileInfo "".path type.string "".ctxt   type.*"".Context p�opDo � �>HE  `� Tgclocals·6d46c0650eba7dbebc0db316e0e0cf3b Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�,"".(*Context).openFile  �  �dH�%    H;a�-  H��HH�T$XH�L$`1�H�\$hH�\$p1�H�\$xH��$�   H�\$PH���   1�H9�tAH�$H�L$H�H����H�l$H�T$H�L$ H�D$(H�l$hH�T$pH�L$xH��$�   H��H�H�$H�L$�    H�L$H�D$H�T$ H�T$@H�D$8H�� t1�H�\$hH�\$pH�D$xH��$�   H��H�H�L$0H�    1�H9�t#H�\$0H�\$pH�D$h1�H�\$xH��$�   H��H�H�    H�$H�    H�\$H�    H�\$�    H�D$��    ����������
      �       �  os.Open   �  <go.itab.*os.File.io.ReadCloser   �  type.*os.File   �  $type.io.ReadCloser   �  <go.itab.*os.File.io.ReadCloser   �   runtime.typ2Itab   �  0runtime.morestack_noctxt   p�  "".autotmp_0039 /type.*os.File "".err type.error "".~r2 Ptype.error "".~r1 0$type.io.ReadCloser "".path type.string "".ctxt   type.*"".Context 6�x��J��5��/� � $�<A"e  ^� Tgclocals·5cbd57cf8f9b35eac9551b20a42afe1f Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60   :$GOROOT/src/go/build/build.go�("".(*Context).isFile  �  �dH�%    H;avrH��XH�\$`H�$H�\$hH�\$H�\$pH�\$�    H�T$H�L$ H�D$(H�\$0H�\$PH�D$HH�� t
�D$x H��X�H�L$@H�$H�T$8H�Z ���D$xH��X��    �u��������
      b  ,"".(*Context).openFile   �       �  0runtime.morestack_noctxt   @�  
"".err type.error "".f ?$type.io.ReadCloser "".~r1 0type.bool "".path type.string "".ctxt   type.*"".Context �O��� �  �;

 
 0` Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�("".(*Context).gopath  �  �dH�%    H�D$�H;A�:  H���   H��$�   1�H��$�   H��$�   H��$   1�H��$�   H��$�   H��$�   H�$H�� ��  H�X0H�|$H�H�H�KH�O�    H�L$H�D$ H�T$(H��$�   H��$�   H��$�   H��$�   H�D$H    H��$�   H�D$@H��$�   H�L$PH�\$HH�l$@H9���   H�\$PH�� �K  H�L�KH�L$xI�� tjH��$�   H�� �   H�K H�C(I9���   H�l$xH�,$L��$�   L�L$H��$�   H�L$H��$�   H�D$�    L��$�   �\$ �� tfH�\$PH��H�\$PH�\$HH��H�\$HH�\$HH�l$@H9��G���H��$�   H��$�   H��$�   H��$�   H��$�   H��$   H���   �L�D$xL�D$XL��$�   H�=    H�|$hH��   L�L$`H�D$pI9��#  L9��  H9��  L��$�   L�$H��$�   H�D$H�|$H�D$�    L��$�   �\$ H��< ����H��$�   H��$�   H��$�   H��H��H9�wBH��$�   H��H��Hk�H�L�KH�l$x�=     uH�+����H�$H�l$�    ����H�-    H�,$H�L$H�D$H�T$H�\$ �    L��$�   H�L$(H�D$0H�T$8H��H��H��$�   H��$�   H��$�   �h���1��.����    1�� ��������������� �����    ��������
      �  6"".(*Context).splitPathList   �   runtime.eqstring   �  go.string."~"   �	   runtime.eqstring   �
 (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0052  type.string "".autotmp_0051 �type.string "".autotmp_0050 �type.*string "".autotmp_0049 �type.int "".autotmp_0048 �type.int "".autotmp_0047  type.string "".autotmp_0043 �type.[]string "".autotmp_0042 _type.[]string "strings.prefix·3 �type.string strings.s·2 �type.string "".p �type.string "".all /type.[]string "".~r0 type.[]string "".ctxt   type.*"".Context "������ � H�A�p.28!�M-.-.^   ���)F1 Tgclocals·087344e727b14a841dc6a2833d52f059 Tgclocals·e2234b98cb6fbb40cb1b6c335fab0a3e   :$GOROOT/src/go/build/build.go�*"".(*Context).SrcDirs  �  �dH�%    H�D$�H;A��  H���   1�H��$  H��$  H��$  1�H��$�   H��$�   H��$�   H��$   H�[(H�� �e  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$�      HǄ$�      H��$   H�� �(  H�k H��$�   H�D$H�l$H�-    H�,$�    H��$   H�$H��$�   H�\$H��$�   H�\$H��$�   H�\$�    H�L$ H�D$(H��$   H�$H�L$xH�L$H��$�   H�D$�    �\$�� ��  H��$�   H��$�   H��$�   H��H��H9��  H��$�   H��H��Hk�H�H��$�   H�kH�l$x�=     ��  H�+H��$   H�$�    H�D$H�l$H�L$H��$�   H��$�   H��$�   H��$�   1�H��$�   H�l$@H��$�   H�l$@H9���  H�D$PH�� �D  H�H�hH�L$HH��$�   H�T$XH��$�   H�l$`H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$�      HǄ$�      H��$�   H�l$`H�hH�l$X�=     ��  H�(H��$   H�$H�D$H��$�   H�\$H��$�   H�\$�    H�L$ H�D$(H��$   H�$H�L$hH�L$H�D$pH�D$�    �\$�� �  H��$�   H��$�   H��$�   H��H��H9���   H��$�   H��H��Hk�H�H�l$pH�kH�l$h�=     uZH�+H�D$PH�L$HH��H��H�l$@H9��k���H��$�   H��$  H��$�   H��$  H��$�   H��$  H���   �H�$H�l$�    �H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�D$0H�T$8H��H��H��$�   H��$�   H��$�   �����>���H�$H�l$�    H��$�   �`���� ����H�$H�l$�    �.���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�D$0H�T$8H��H��H��$�   H��$�   H��$�   ����������������    ���������>
      �  type.[2]string   �  "runtime.newobject   �  """.statictmp_0062   � """.statictmp_0062   �  """.statictmp_0062   �0 """.statictmp_0062   �  type.string   �  (runtime.typedmemmove   �  ,"".(*Context).joinPath   �  &"".(*Context).isDir   � (runtime.writeBarrier   �  ("".(*Context).gopath   �	  type.[2]string   �	  "runtime.newobject   �
  """.statictmp_0069   �
 """.statictmp_0069   �
  """.statictmp_0069   �
0 """.statictmp_0069   � (runtime.writeBarrier   �  ,"".(*Context).joinPath   �  &"".(*Context).isDir   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  0runtime.morestack_noctxt   @�   "".autotmp_0070  type.*[2]string "".autotmp_0068 �type.[]string "".autotmp_0067 �type.string "".autotmp_0066 �type.*string "".autotmp_0065 �type.int "".autotmp_0064 �type.int "".autotmp_0061 �type.[]string "".autotmp_0060  type.bool "".autotmp_0059 _type.[]string "".autotmp_0058  type.[]string "".dir �type.string "".p �type.string "".dir �type.string "".all /type.[]string "".~r0 type.[]string "".ctxt   type.*"".Context "������ �
 j�9�6]��3V8VV	 B t�82|��/�&E"	)Q Tgclocals·cffcb3fa139580cffca8ac28af4ff263 Tgclocals·605a1b837cd4aeeb8235060aa13f27b7   :$GOROOT/src/go/build/build.go�""".defaultContext  �  �dH�%    H��$���H;A�*  H��p  H��$x  W�H����    H��$�   W�H����    H�    H�$H�D$   H�    H�\$H�D$   �    H�L$ H�D$(H��$�   H��$�   H�    H�$H�D$   H�    H�\$H�D$   �    H�L$ H�D$(H��$�   H��$�   �    H�$H�D$H�L$xH�$H��$�   H�D$�    H�L$H�D$H��$�   H��$�   H�    H�$H�D$   1�H�\$H�\$�    H�L$ H�D$(H��$�   H��$�   H�    H��$�   HǄ$�      H�    H�$�    H�|$H��H�� ��  H�5    �    H�� ��  H��   H��   H��$�   H��$  H��$�   H��$  H��$�   H��$   H�    H�$H�D$   �    H�L$H�D$H�L$xH�L$hH��$�   H��ubH�l$hH�,$H�D$pH�D$H�-    H�l$H�D$   �    H�D$p�\$ �� t&1ۈ�$�   H��$�   H��$x  �    H��p  �H��uGH�l$hH�,$H�D$pH�D$H�-    H�l$H�D$   �    �\$ �� tH��   ��$�   �H��$�   H��$�   H���8  H�-    H�,$H�D$   H�L$hH�L$H�D$pH�D$�    �\$ �� ��   H��$�   H��$�   H����   H�-    H�,$H�D$   H�L$hH�L$H�D$pH�D$�    �\$ �� ��   H�\$HH�$H��$�   H�|$H�H�H�KH�OH�    H�\$H�D$    H��$�   H�|$(H�H�H�KH�O�    H�L$8H�D$@H�    H�$H�    H�\$H�L$hH�L$H�D$pH�D$�    H�\$ �+@��$�   �D���1ۈ�$�   �6�����q�����T����    �����F
      d�  runtime.duffzero   ��  runtime.duffzero   �  $go.string."GOARCH"   �  "go.string."amd64"   �  "".envOr   �   go.string."GOOS"   �  "go.string."linux"   �  "".envOr   �  runtime.GOROOT   �  path.Clean   �  $go.string."GOPATH"   �  "".envOr   �  go.string."gc"   �  type.[6]string   �  "runtime.newobject   �  """.statictmp_0086   ��  runtime.duffcopy   �  .go.string."CGO_ENABLED"   �  os.Getenv   �  go.string."0"   �	   runtime.eqstring   �	�  runtime.duffcopy   �
  go.string."1"   �
   runtime.eqstring   �  "go.string."amd64"   �   runtime.eqstring   �  "go.string."linux"   �   runtime.eqstring   �  go.string."/"   �  *runtime.concatstring3   �  (type.map[string]bool   �  "".cgoEnabled   �  4runtime.mapaccess1_faststr   �  0runtime.morestack_noctxt   ��  "".autotmp_0091 �type.[32]uint8 "".autotmp_0090  type.string "".autotmp_0089  type.string "".autotmp_0088  type.string "".autotmp_0085 �type.[]string "".autotmp_0083  type.string "".autotmp_0082  type.string "".autotmp_0081  type.string "".autotmp_0080 �type.string "".autotmp_0079  type.string "".autotmp_0078  type.string "".autotmp_0077 �type.string "".c �type."".Context "".~r0  type."".Context ""������ � `�6HHC?v5B	=��	  s�h� Tgclocals·7353ec067a80b85e773ae30131808ed8 Tgclocals·b747f90b0df18c3781c6f6b1a3b90488   :$GOROOT/src/go/build/build.go�"".envOr  �  �dH�%    H;av`H�� 1�H�\$HH�\$PH�\$(H�$H�\$0H�\$�    H�L$H�D$H�� uH�\$8H�\$HH�\$@H�\$PH�� �H�L$HH�D$PH�� ��    �����������
      f  os.Getenv   �  0runtime.morestack_noctxt   `@  "".~r2 @type.string "".def  type.string "".name  type.string @L?@? � �"	 
 2N Tgclocals·b4c25e9b09fd0cf9bb429dcefe91c353 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�."".(*Package).IsCommand  �  �dH�%    H;avcH��8H�\$@H�� tPH�KH�kH��u;H�L$(H�$H�l$0H�l$H�    H�\$H�D$   �    �\$ �\$HH��8��D$H ����    ��������
      �   go.string."main"   �   runtime.eqstring   �  0runtime.morestack_noctxt    p  "".autotmp_0092 type.string "".~r0 type.bool "".p   type.*"".Package pSopo � �_ 
 T, Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad   :$GOROOT/src/go/build/build.go�."".(*Context).ImportDir  �  �dH�%    H;avzH��H1�H�\$xH��$�   H�\$PH�$H�    H�\$H�D$   H�\$XH�\$H�\$`H�\$ H�\$hH�\$(�    H�T$0H�L$8H�D$@H�T$pH�L$xH��$�   H��H��    �m����������������
      \  go.string."."   �  ("".(*Context).Import   �  0runtime.morestack_noctxt   p�  
"".~r3 Ptype.error "".~r2 @ type.*"".Package "".mode 0$type."".ImportMode "".dir type.string "".ctxt   type.*"".Context �u� � �"g 
 ^B Tgclocals·b60dc0a6046c556b02baa766a3fd5a27 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�*"".(*NoGoError).Error  �  �dH�%    H;avcH��81�H�\$HH�\$PH�$    H�    H�\$H�D$    H�t$@H�|$H�H�H�NH�O�    H�\$(H�\$HH�\$0H�\$PH��8��    ��������
      T  Xgo.string."no buildable Go source files in "   �  *runtime.concatstring2   �  0runtime.morestack_noctxt   0p  "".~r0 type.string "".e  $type.*"".NoGoError p^o � �S 
 T, Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�@"".(*MultiplePackageError).Error  �  �dH�%    H�D$�H;A��  H���   1�H��$�   H��$�   H�|$xW�H����    H�\$xH�� ��  H�D$h   H�D$p   H�\$`H�    H�$H��$�   H�� �j  H�KH�CH�k H�l$XH�L$HH�� H�D$P�>  H�L$H�D$    �    H�L$H�D$ H�\$`H�L$8H�H�D$@�=     ��  H�CH�    H�$H��$�   H�� ��  H�K(H�C0H�k8H�l$XH�L$HH�� H�D$P��  H�L$H�D$    �    H�L$H�D$ H�\$`H��H�L$8H�H�D$@�=     �@  H�CH�    H�$H��$�   H�� �  H�KH�CH�k H�l$XH��H�L$HH��H�D$P��  H��H�\$H�D$    �    H�L$H�D$ H�\$`H�� H�L$8H�H�D$@�=     ��  H�CH�    H�$H��$�   H�� �f  H�K(H�C0H�k8H�l$XH��H�L$HH��H�D$P�7  H��H�\$H�D$    �    H�L$H�D$ H�\$`H��0H�L$8H�H�D$@�=     ��   H�CH�    H�$H��$�   H�\$H�|$ ��   H�D$    �    H�L$H�D$ H�\$`H��@H�L$8H�H�D$@�=     u]H�CH�    H�$H�D$(   H�\$`H�\$H�\$hH�\$H�\$pH�\$ �    H�L$(H�D$0H��$�   H��$�   H���   �L�CL�$H�D$�    듉%    �L���L�CL�$H�D$�    �����    �����L�CL�$H�D$�    �_����    ������L�CL�$H�D$�    �����    ��6���L�CL�$H�D$�    �����    �������T����    ��������������:
      |�  runtime.duffzero   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �	  runtime.convT2E   �	 (runtime.writeBarrier   �
  type.string   �
  runtime.convT2E   � (runtime.writeBarrier   �  hgo.string."found packages %s (%s) and %s (%s) in %s"   �  fmt.Sprintf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0�  "".autotmp_0104  "type.interface {} "".autotmp_0103  "type.interface {} "".autotmp_0102  "type.interface {} "".autotmp_0101  "type.interface {} "".autotmp_0100 �"type.interface {} "".autotmp_0099 �(type.[5]interface {} "".autotmp_0096 �&type.[]interface {} "".~r0 type.string "".e  :type.*"".MultiplePackageError "������ � �1� 2 ��4*


( Tgclocals·cb395d89503762333b1bfb09ba74eb12 Tgclocals·345f1bd1394e1f5bdb891635a73ee227   :$GOROOT/src/go/build/build.go�"".nameExt  �  �dH�%    H;a��   H��(1�H�\$@H�\$HH�\$0H�$H�\$8H�\$H�    H�\$H�D$   �    H�D$ H�� }1�H�\$@H�\$HH��(�H�l$8H9�w!L�D$0H)�H�� tM� L�D$@H�l$HH��(��    �    �X�����������

      r  go.string."."   �  "strings.LastIndex   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @P  "".~r1  type.string "".name  type.string PTOP*OPO � �#22	 
 Ke Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�("".(*Context).Import  ��  ��dH�%    H��$(���H;A��  H��X  W�H��$X	  �    G�H��$x  �    G��$p  �$0  �$@  1�H��$�  H��$�  H�    H�$�    H�|$H��H�� ��  W��    G�H��$�  H��$p  H�hHH��$h  �=     �H  H�h@H��$  H��$p  H�� �L  H��$h  H��$�  H��$p  H��$�  1�H��$p  H��$x  H��$p  H�� �  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     uvH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$  H��$�  H��$�  H��$�  H��X  �L�CL�$H�D$�    �w���������1�H��$   H��$(  1�H��$@  H��$H  1�H��$0  H��$8  1�H��$P  H��$X  H��$`  H���   H�� tlH��$h  H�$H�    H�\$H�D$   H��$`  H�� �G}  H���   H�|$H�H�H�KH�O�    H�\$(H��$P  H�\$0H��$X  H��$`  H�� ��|  H�KHH��$P  H�CPH���z  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$`  H��$P  H��$X  �\$ �� ��y  H�$    H�    H�\$H�D$   H�� ��y  H�ZH�|$H�H�H�KH�OH�    H�\$(H�D$0   H�|$8H�
H�H�JH�OH��$P  H�\$HH��$X  H�\$P�    H�T$XH�L$`1�H��$X	  H��$`	  H��$h	  H��$p	  H��$x	  H��$�	  H��$X	  H�-    H�(H��$`  H�hH��$  H�hH��$@  H�hH��$   H�P H��$(  H�H(H��$�  H�H����Ƅ$�    L��$h  L��$p  H��$p  H��$x  H���^x  L�$H�L$H�    H�\$H�D$   �    L��$p  H��$x  �\$ H��< �x  H����w  L�$H�L$H�    H�\$H�D$   �    L��$p  H��$x  �\$ H��< ��w  L��$   H�=    H��$   H��   H��$(  H��$  H9��qw  H9��aw  H9��Qw  L��$P  L�$H��$X  H�D$H�|$H�D$�    L��$p  H��$x  �\$ H��< ��v  L��$�  H�5    H��$�  H��   H��$�  H��$�  H9���v  H9���v  H9���v  L��$P  L�$H��$X  H�D$H�t$H�D$�    �\$ H��< ��]  1�H��$@  H��$H  H��$�  H�� �L  H��$h  H��$�  H��$p  H��$�  1�H��$p  H��$x  H��$p  H�� �  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     uvH�CH�    H�$H�D$/   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$  H��$�  H��$�  H��$�  H��X  �L�CL�$H�D$�    �w���������H��$`  H�$H��$h  H�\$H��$p  H�\$�    �\$�� �1\  H�    H�$�    H�D$H�� �\  HǄ$x     HǄ$�     H��$p  H��$�  H�hH��$x  �=     ��[  H�(H��$p  H��H��H�kH��$h  �=     �i[  H�+H��$`  H�$H�D$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� �[  H��$X  H�CH��$P  �=     ��Z  H�H�    H��$  H��$`  H�[(H�� ��S  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$x     HǄ$�     H��$`  H�� �FZ  H�k H��$p  H�D$H�l$H�-    H�,$�    H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$`  H�$H��$�  H�L$H��$�  H�D$H��$  H�|$H�H�H�NH�O�    H�T$(H��$`  H�L$0H��$h  �\$8�� �CR  H�$H�L$H��$  H���H��$  �\$�� �R  H��   @���   H��$h  H�iHH��$`  �=     ��Q  H�i@H��$`  H�� ��Q  H�k H�� ��Q  L�APL�D$H�l$H�-    H�,$�    H��$  H�[XH�� �o  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$x     HǄ$�     H��$  H�� ��P  H�kPH��$p  H�D$H�l$H�-    H�,$�    H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� �qP  H��$X  H�ChH��$P  �=     �9P  H�K`H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$x     HǄ$�     H��$  H�� ��O  H�kPH��$p  H�D$H�l$H�-    H�,$�    H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� �CO  H��$X  H�CxH��$P  �=     �O  H�KpH�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$x     HǄ$�     H��$  H�� ��N  H�kPH��$p  H�D$H�l$H�-    H�,$�    H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� �N  H��$X  H���   H��$P  �=     ��M  H���   H��$H  H�� �<  H�    H�$�    H�D$H�� ��M  HǄ$x     HǄ$�     H��$  H�� �gM  H�kPH��$p  H�D$H�l$H�-    H�,$�    H��$p  H��$(  H��H�kH��$   �=     �M  H�+H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� ��L  H��$X  H���   H��$P  �=     �eL  H���   H�    H�$�    H�D$H�� �8L  HǄ$x     HǄ$�     H��$  H�� �L  H�kPH��$p  H�D$H�l$H�-    H�,$�    H��$p  H��$H  H��H�kH��$@  �=     ��K  H�+H��$`  H�$H��$p  H�\$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$  H�� �CK  H��$X  H���   H��$P  �=     �K  H���   H��$�  H��H�� t8H��$  H��$�  H��$0  H��$�  H��$8  H��$�  H��X  À�$�    tJH��$�  H��H�� t8H��$  H��$�  H��$0  H��$�  H��$8  H��$�  H��X  �H��$`  H�$H��$  H�|$H�H�H�NH�O�    H�\$H��$  H�\$ H��$  H�\$(H��$   H�\$0H��$  H�\$8H��$  H��$  H�� t8H��$  H��$�  H��$  H��$�  H��$  H��$�  H��X  �1�H��$�  H��$�  1�H��$`  H��$h  H��$p  1�H��$�  H��$�  1�H��$�  H��$�  H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$  H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�  H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�  1�H��$(	  ��$0	  ��$1	  ��$4	  H��$8	  H��$@	  H��$H	  H��$P	  H��$�
  W�H����    G�H�    H�$H�D$    H��$(	  H�\$H��$�
  H�\$�    H�\$ H��$�  HǄ$�      H�    H�$�    H�\$H��$�  H��$�  H�� ��G  W��    H��$�  H�C   H��$�  H��$�  H��$�  H��$�  H��$�  H��$   H��$  H��$  H��$  H��$   H��$   H��$(  H��$   1�H��$`  H��$  H��$�  H��$`  H9���   H��$�  H�� �G  H�+H��$   H�kH��$(  H��$  H��$   H��$�  H��$(  H��$�  H��$�  H�$H��$�  H�[ ���\$�� �	  H��$�  H��H��$�  H��$  H��H��$`  H9��W���H��$�  H�� t8H��$  H��$�  H��$�  H��$�  H��$�  H��$�  H��X  �H��$  H���   H��$  H��   H��$  H���  H��$H  H��$  H���  H��$@  H��$H  H��H�H�H��$@  H�H�� �  H�    H�$�    H�\$H��$P  H��$  H�� ��   H��$P  H�� ��   H�\$H�l$H�-    H�,$�    H��$P  H��$P  H�    H��$p  H��$p  1�H9�t8H��$  H��$�  H��$P  H��$�  H��$p  H��$�  H��X  �H�    H�$H�    H�\$H�    H�\$�    H�\$H��$p  둉�B����E �(���H��$�  H��$�  H��$`
  W�H����    H�    H�$H��$�  H�\$H��$`
  H�\$�    H��$`
  1�H9���   H��$`
  H�� ��  H�+H��$�  H�kH��$�  H��$  H���   H���   H���   H��H��H9���  H���   H��H��Hk�H�H��$�  H�kH��$�  �=     �i  H�+H��$`
  H�$�    H��$`
  1�H9��O���H��$  H�� �)  H���   H�H�$H�KH�L$H�KH�L$�    H��$  H�$�    H�D$H�T$H�L$H�\$ H��$H  H��$  H�� ��  H��$`  H���  H��$h  H���  H��$X  �=     �q  H��x  H��$  H�� �Q  H��$H  �=     �"  H���  H��$�  H�$�    H�D$H�T$H�L$H�\$ H��$H  H��$  H�� ��  H��$`  H���  H��$h  H���  H��$X  �=     ��  H���  H��$  H�� �h  H��$H  �=     �9  H���  H��$�  H�$�    H��$  H�D$H�T$H�L$H�\$ H��$H  H�� ��  H��$`  H���  H��$h  H���  H��$X  �=     ��  H���  H�� �  H��$H  �=     �H  H��   H��   H��$@  H��$@  H�� ��  H���  H���  H���  H��$X  H��H��$`  H��$h  H��H��$x  H��$h  H�H)�H�� ~SH�    H�$H��$p  H�t$H�T$H��$�  H�L$H�D$ �    H��$`  H�t$(H�\$0H��$x  H�L$8H�    H�$L��$h  H��H��L�I��H��$�  H9��G  H9��>  H)�I)�I��H��$p  I�� tHk�I�H�l$L�D$L�L$H��$`  H�\$ H��$h  H�\$(H��$p  H�\$0�    H��$�  H��$`  H��$h  H�H9���   H��H��$  H���  H���  H��$p  �=     uvH���  H��$  H�� t]H���  H�H�$H�KH�L$H�KH�L$�    H��$  H��$�  H��$0  H��$�  H��$8  H��$�  H��X  É�L���  L�$H�l$�    �w����    �    L��   L�$H�l$�    H��$  ������z���L���  L�$H�D$�    H��$  �N��������L���  L�$H�l$�    ���������L���  L�$H�D$�    �e�����$���L���  L�$H�l$�    ����������L��x  L�$H�D$�    �|�����;���������H�$H�l$�    ����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���   H���   H��$@  �=     uH���   �����L���   L�$H�T$�    H��$@  H��$�   �����뙉�]���H��$�  H�$H��$�  H�[8��H�\$H��$�  H�\$H��$�  H��$�  H�$H��$�  H�\$�    H��$  H�\$H��$�  H�\$H��$�  1�H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H�-    H�+H��$�  H��$�  H�kH��$�  H�CH��$�  H��$�  H�kH��$�  H�k H��$�  H��$8  H��$`  H�$H�|$H�H�H�HH�OH��$�  H�\$H��$�  H�\$ �D$(H��$�  H�\$0�    �\$8��$�   H�\$@H��$(  H�\$HH��$0  H�\$PH��$8  H�\$XH��$�  H�\$`H��$�  H�\$hH��$   H�\$pH��$(  H��$   H�� t+H��$   H�$H��$(  H�\$H��$8  H����������$�    �o  H��$�  H�������H��$�  H�,$H��$�  H�l$H�-    H�l$H�D$   �    �\$ �� �����H��$  H��  H��  H��   H��H��H9�wLH��  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�9���H�$H�l$�    �&���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��  H��   H��$@  �=     uH��  �A���L��  L�$H�T$�    H��$@  H��$�   ������H��$�  H��$P  H��$�  H��|TH����3  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  H�\$ H�� ��3  H��|TH����.  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  H�\$ H�� �n.  H���  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� ��   H��$`  H��$h  H��$p  H��H��H9�wMH��$h  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+����H�$H�l$�    �����H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$h  H��$p  H��$`  �e���H���e  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �  H��$  H��@  H��H  H��P  H��H��H9�wLH��H  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��H  H��P  H��$@  �=     uH��@  �A���L��@  L�$H�T$�    H��$@  H��$�   ������H��$X  H���M  H�$H�D$H�-    H�l$H�D$   �    �\$ �� �  H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+����H�$H�l$�    �s���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   ������H��$(  H��$   H��$0  H��$  H��$8  H��$  H�    H�$H��$   H�\$H�D$    �    H�\$H�|$H�H�H�KH�OH��$   H�$H��$�  H�\$H��$�  H�\$H�D$(   �    H�\$0H��$   H�\$8H��$   H�\$@H��$(  H��$   H�� t+H��$   H�$H��$(  H�\$H��$8  H��������H��$   H�kH�� �g)  H�]H��$P  H�]H��$X  H��$X  H���]  H��$P  H�,$H��$X  H�l$H�-    H�l$H�D$   �    �\$ �� �  H��$  H��  H��  H��   H��H��H9�wLH��  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��  H��   H��$@  �=     uH��  �A���L��  L�$H�T$�    H��$@  H��$�   ������H��$�  H��$�  H��$�  H��$�  H�    H��$0  HǄ$8     �D$| H��$�  H��$8  H9���'  H��$�  H��$H  H��$8  H��$@  H��$H  H��$@  H)�H��$8  H��$8  H��$�  H9��%'  L��$�  H)�H�� tM�H��H��H��$8  H9���&  L��$P  L�$H��$X  H�D$H��$0  H�\$H��$8  H�\$�    �\$ H�؈D$|�\$|��$�   Ƅ$�    ��$�    �c  H��$P  H��$  H��$X  H��$  H�    H��$@  HǄ$H     �D$} H��$  H��$H  H9��,&  H��$  H��$0  H��$H  H��$(  H��$0  H��$(  H)�H��$   H��$   H��$  H9���%  L��$  H)�H�� tM�H��$�  L��$�  H��$�  H��$H  H9���%  H��$�  H�$H��$�  H�\$H��$@  H�\$H��$H  H�\$�    �\$ H�؈D$}�|$} t-Ƅ$�   H��$X  H��$X  H��H9��%  H��$X  H��$  H�[H�� �    H��$  H��$X  H�kH��$P  �=     ��  H�kH��$�  H��$�  H��$�  H��$�  H��$   H�] 1�H9���   H��$  H�[8H�� ��   H��$   H�+H�,$�    H�\$H��$  H�\$H��$  H��$  H�$H��$  H�\$�    H�\$H��$�  H�\$H��$�  H��$  H��$�  H�k8H��$�  �=     ��  H�k0H��$�  H��H�� �x  H��$(  H�$H��$0  H�\$H��$8  H�\$�    H�\$H��$�  H�\$ H��$�  H�\$(H��$�   H��$�   H�� �  H��$�  H�$H��$�  H�\$�    H�\$H��$�  H�\$H��$�  H�\$ H��$�  H�\$(H��$�  H��$�  H�� �T  H��$�  H��$�  H��$�  H��$�  H��$�   H��$  1�H��$�  H��$�  H��$�  H��$�  H��$�  H�� ��  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     �Z  H�CH�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$`  H�H��$h  �=     ��  H�CH�    H�$H�D$"   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$�  H�$H��$�  H�D$H��$8  H���Ƅ$�    H��$   H�� �N  H�kH��$�  H�k H��$�  H�k(H��$�  HǄ$X      H��$�  H��$P  H��$�  H��$`  H��$X  H��$P  H9���   H��$`  H�� ��  H�+H��$   H�kH��$  H��$   H��$�  H��$  H��$�  HǄ$�      H��$�  1�H9�tH�[H�-    H9��P  H��$�  H��$�  �D$~H��$�  H��$(  �|$~ �e  H��$`  H��H��$`  H��$X  H��H��$X  H��$X  H��$P  H9�������$�    ��  H�    H��$�  HǄ$�     Ƅ$�   H�    H�$H��$�  H�\$H��$�  H�\$H��$�   H�\$�    H��$`  �]@�� �  H��$  H���   H��   H��  H��H��H9�wLH��   H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+����H�$H�l$�    �}���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��   H��  H��$@  �=     uH���   �A���L���   L�$H�T$�    H��$@  H��$�   ������H��$  H��  H��  H��   H��H��H9�wLH��  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�t���H�$H�l$�    �a���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��  H��   H��$@  �=     uH��  �A���L��  L�$H�T$�    H��$@  H��$�   �����뙀�$�    �  H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�J���H�$H�l$�    �7���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   �����뙀�$�    �  H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+� ���H�$H�l$�    ����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   ������H��$  H���   H���   H���   H��H��H9�wLH���   H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���   H���   H��$@  �=     uH���   �A���L���   L�$H�T$�    H��$@  H��$�   ������H��$(  H�� ��  H�k H��$�  H�k(H��$�  H�k0H��$�  HǄ$       H��$�  H��$�   H��$�  H��$X  H��$   H��$�   H9�� ���H��$X  H�� �   H�+H��$�  H�kH��$�  H��$�  H��$@  H��$�  H��$H  HǄ$�      H��$@  1�H9�tH�[H�-    H9���  H��$H  H��$�  �D$H��$�  H��$�  �|$ u,H��$X  H��H��$X  H��$   H��H��$   ����H��$�  H�kH�� �.  H�]H��$�  H�]H��$�  H��$�  H�$H��$�  H�\$�    H�\$H��$`  H�\$H��$h  H�\$ H��$�  H�\$(H��$�  H��$�  H�� ��  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  1�H��$x  H��$�  H��$�  H��$�  H��$x  H�� �7  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     ��  H�CH�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$`  H�H��$h  �=     �1  H�CH�    H�$H�D$/   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    ��$�    ��  H��$`  H��$�  H��$h  H��$�  H��$`  H��$�  H��$h  H��$�  H�    H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H�� �6  H�+H��$�  H�kH��$�  H�kH��$�  H��$�  H��$�  HǄ$�       H��$�  H�]1�H9���  H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   H��$   H�$H��$�   H�\$�    H�\$H��$ 	  H�\$H��$	  H�\$ H��$	  H�\$(H��$	  H�\$0H��$ 	  H��$�  H��$�  H��$�  H��H��H9��w  H��H��H��$�  H��$�  H��$�  H��H��Hk�(H�H��$	  H�kH��$	  H�kH��$	  H�kH��$ 	  H�k H��$ 	  �=     ��  H�+H�    H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H��$h  H���3���H��$`  H�,$H��$h  H�l$H�-    H�l$H�D$   �    �\$ �� �������$�    �O  H��$�  H��$�  H��$�  H��$�  1�H��$0  H��$8  H��$0  H�� �  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     uyH�CH�    H�$H�D$#   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$�  H�$H��$�  H�D$H��$8  H�������L�CL�$H�D$�    �t���������H��$�  H�+H��$0  H��$0  1�H9�u5H��$(  H�k(H��$  H��$  H��uH��$(  H�+H��$0  H��$0  1�H9���   H��$`  H�$H��$�  H�\$H��$�  H�\$H��$  H�\$H��$0  H�\$ �    H�\$(H��$   H�\$0H��$  H��$   H�� t&H��$   H�$H��$  H�\$H��$8  H���Ƅ$�   ����H�$H�l$�    �����H�-    H�,$H�T$H�D$H�L$H�\$ �    H�T$(H�D$0H�L$8�Q���H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   �s�����������$�    �  H��$`  H��$�  H��$h  H��$�  H��$`  H��$�  H��$h  H��$�  H�    H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H�� �z  H�+H��$�  H�kH��$�  H�kH��$�  H��$�  H��$�  HǄ$�       H��$�  H�]1�H9���  H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   H��$   H�$H��$�   H�\$�    H�\$H��$ 	  H�\$H��$	  H�\$ H��$	  H�\$(H��$	  H�\$0H��$ 	  H��$�  H��$�  H��$�  H��H��H9���   H��H��H��$�  H��$�  H��$�  H��H��Hk�(H�H��$	  H�kH��$	  H�kH��$	  H�kH��$ 	  H�k H��$ 	  �=     u?H�+H�    H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    �.���H�$H�l$�    �H�-    H�,$H�T$H�D$H�L$H�\$ �    H�T$(H�D$0H�L$8����H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   �/��������H��$`  H��$�  H��$h  H��$�  H��$`  H��$�  H��$h  H��$�  H�    H�$H��$  H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H�� �z  H�+H��$�  H�kH��$�  H�kH��$�  H��$�  H��$�  HǄ$�       H��$�  H�]1�H9���  H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   H��$   H�$H��$�   H�\$�    H�\$H��$ 	  H�\$H��$	  H�\$ H��$	  H�\$(H��$	  H�\$0H��$ 	  H��$�  H��$�  H��$�  H��H��H9���   H��H��H��$�  H��$�  H��$�  H��H��Hk�(H�H��$	  H�kH��$	  H�kH��$	  H�kH��$ 	  H�k H��$ 	  �=     u?H�+H�    H�$H��$  H�\$H��$�  H�\$H��$�  H�\$�    �'���H�$H�l$�    �H�-    H�,$H�T$H�D$H�L$H�\$ �    H�T$(H�D$0H�L$8����H��$�  H�kH��$�  HǄ$�       H��$�  H�+H��$�   H��$�   H��$�   H��$�   H��$�   �/��������L�CL�$H�D$�    ����L�CL�$H�D$�    �E����������E �����HǄ$�      �D$ �[�����������W���HǄ$�      �D$~ ������-��������L�CL�$H�D$�    �
���L�CL�$H�D$�    ���������H��$  H�[(H�� ubH��$  H��$�  H�k(H��$�  �=     u)H�k H��$�  H��$�  H��$�  H��$�  �����L�C L�$H�l$�    ��H��$  H�� �&  H�k H��$�  H�k(H��$�  H��$�  H��$�  H9�uFH��$�  H�,$H��$�  H�l$H��$�  H�l$H��$�  H�l$�    �\$ �� �c���H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$
  W�H����    H��$
  H��$h  H��$h  H�� �  HǄ$�     HǄ$�     H��$�  H�    H�$H��$  H�\$H�|$ ��  H�D$ H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     �i  H�CH�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$`  H�H��$h  �=     ��  H�CH�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H�� H��$`  H�H��$h  �=     �{  H�CH�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��0H��$`  H�H��$h  �=     �  H�CH�    H�$H��$  H�\$H�|$ ��   H�D$    �    H�L$H�D$ H��$�  H��@H��$`  H�H��$h  �=     uyH�CH�    H�$H�D$/   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$�  H�$H��$�  H�D$H��$8  H����B���L�CL�$H�D$�    �t����%    �$���L�CL�$H�D$�    �����L�CL�$H�D$�    �r���L�CL�$H�D$�    �����L�CL�$H�D$�    �����%    �.���������������L�C0L�$H�l$�    ����L�CL�$H�l$�    ����H��$  H�� ��  H�kH��$  H�kH��$  H��$X  H��$  H9�uFH��$P  H�,$H��$X  H�l$H��$  H�l$H��$  H�l$�    �\$ �� �����H�    H�$�    H�\$H��$x  H��$  H�� �  H��$x  H�� ��  H�\$H�l$H�-    H�,$�    H�    H�$�    H�D$H�� ��  HǄ$x     HǄ$�     H��$  H�� ��  H�kH��$p  H�D$H�l$H�-    H�,$�    H��$p  H��$X  H��H�kH��$P  �=     �$  H�+H��$x  H��$x  H�kH��$�  H�k H��$p  �=     ��  H�kH�    H�$�    H�D$H�� ��  HǄ$x     HǄ$�     H��$p  H��$�  H�hH��$�  �=     �O  H�(H��$�  H��H��H�kH��$�  �=     �	  H�+H��$x  H��$x  H�k0H��$�  H�k8�=     ��  H�C(H��$x  H��$x  H�    H��$p  H��$p  1�H9��R  H��$x  H��$p  H��$�  H�$H��$�  H�D$H��$8  H���H��$  H��(  H��0  H��8  H��H��H9�wLH��0  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��0  H��8  H��$@  �=     uH��(  �A���L��(  L�$H�T$�    H��$@  H��$�   ������H�    H�$H�    H�\$H�    H�\$�    H�\$H��$p  �t���L�C(L�$H�D$�    �+���H�$H�l$�    H��$p  �����H�$H�l$�    H��$p  ����� �N���L�CL�$H�l$�    ����H�$H�l$�    �������o���� �>����������E �������;����    1������    1�����1��G����    1��9����E ����H��|TH���  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  H�\$ H�� ��  H���e  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �  H��$  H��p  H��x  H���  H��H��H9�wLH��x  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�6���H�$H�l$�    �#���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��x  H���  H��$@  �=     uH��p  �A���L��p  L�$H�T$�    H��$@  H��$�   ������H��$X  H�������H�$H�D$H�-    H�l$H�D$   �    �\$ �� �m���H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   ������H���e  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �  H��$  H��X  H��`  H��h  H��H��H9�wLH��`  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�h���H�$H�l$�    �U���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H��`  H��h  H��$@  �=     uH��X  �A���L��X  L�$H�T$�    H��$@  H��$�   ������H��$X  H�������H�$H�D$H�-    H�l$H�D$   �    �\$ �� ���������H��|TH���0  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  H�\$ H�� ��   H��uIH�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �����H��uIH�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �����H��$X  H�������H�$H�D$H�-    H�l$H�D$   �    �\$ �� �C����Z���H��|TH����  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  H�\$ H�� ��  H��uIH�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �����H��$X  H�������H�$H�D$H�-    H�l$H�D$   �    �\$ �� �n���H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�ؼ��H�$H�l$�    �ż��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   ������H���e  H�$H��$X  H�D$H�-    H�l$H�D$   �    H��$P  H��$X  �\$ �� �  H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�i���H�$H�l$�    �V���H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   ������H��$X  H�������H�$H�D$H�-    H�l$H�D$   �    �\$ �� �����H��$  H���  H���  H���  H��H��H9�wLH���  H��H��Hk�H�H��$�  H�kH��$�  �=     uH�+�
���H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$  H�� tcH��H��$�   H��H���  H���  H��$@  �=     uH���  �A���L���  L�$H�T$�    H��$@  H��$�   �����뙉���������L���   L�$H�L$�    �����鶴��H�$H�l$�    �O��������� �����L���   L�$H�L$�    鈳����V���H�$H�l$�    �����钲��� �a���L���   L�$H�L$�    �����������c���L�CpL�$H�L$�    �����鶰����5���L�C`L�$H�L$�    鴯���鈯���������b�����M���L�A@L�$H�l$�    H��$  ����H��$`  H�$�    H�T$H�L$H�D$H��$H  H��$P  H��$X  H��$�  1�H��$x  H��$X  H��$p  H��H��$X  H9�����H��$�  H�� ��  H�H�iH��$`  H��$�   H��$P  H��$�  H��$X  H��$�  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$`     HǄ$h     H��$X  H��$�  H�hH��$�  �=     ��  H�(H��$`  H�$H�D$H��$`  H�\$H��$h  H�\$�    H�L$ H�D$(H��$`  H�$H��$�  H�L$H��$�  H�D$H��$  H�|$H�H�H�NH�O�    H�T$(H��$p  H�L$0H��$x  �\$8�� �  H�$H�L$H��$  H����\$�� ��  H��$`  H�[(H�� ��  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hH�-    H�h H�-    H�h(HǄ$`     HǄ$h     H��$`  H�� �K  H�k H��$X  H�D$H�l$H�-    H�,$�    H��$X  H��$x  H�� H�kH��$p  �=     ��  H�+H��$`  H�$H��$X  H�\$H��$`  H�\$H��$h  H�\$�    H�L$ H�D$(H��$`  H�$H��$�  H�L$H��$�  H�D$�    �\$�� tNH��$  H��$�  H���   H��$�  �=     uH���   鼪��L���   L�$H�l$�    颪��H��$�   H��$X  H9���  H��$H  H��$X  H��$`  H��$h  H��$@  1�H��$8  H��$  H��$0  H��$  H9���  H��$�  H�� ��  H�H�hH��$P  H��$P  H��$0  H��$X  H��$8  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hH�-    H�h H�-    H�h(HǄ$H     HǄ$P     H��$@  H��$8  H�hH��$0  �=     ��  H�(H��$x  H��H�� H�kH��$p  �=     �j  H�+H��$`  H�$H�D$H��$H  H�\$H��$P  H�\$�    H�L$ H�D$(H��$`  H�$H��$�  H�L$H��$�  H�D$�    �\$�� tNH��$  H��$�  H���   H��$�  �=     uH���   鍨��L���   L�$H�l$�    �s���H��$�  H��$P  H��H��H��$  H9�����H��$  H��$x  H�kHH��$p  �=     uIH�k@H��$  H��$�  H�kXH��$�  �=     u	H�kP�����L�CPL�$H�l$�    �ݧ��L�C@L�$H�l$�    �H�$H�l$�    H��$@  �~���H�$H�l$�    H��$@  �8���� �h����    H�$H�l$�    ���������H��$�  H��$`  H��H���R���H�$H�l$�    H��$X  ������S����鳥��H�$H�L$�    ���������H�$H�l$�    H��$p  ����H�$H�l$�    H��$p  �9���� �����Ȥ��H��$h  H��$   H��$p  H�5    H��$  H��   H��$  H��$  H9��:  H9��*  H9��  H��$P  H�<$H��$X  H�D$H�t$H�D$�    �\$ H��< �L  H��$h  H��$�  H��$p  H��$�  1�H��$p  H��$x  H��$p  H�� �  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     uvH�CH�    H�$H�D$&   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$  H��$�  H��$�  H��$�  H��X  �L�CL�$H�D$�    �w���������1�H��$�	  H��$�	  H��$�	  H��$�	  H��$�	  H��$�	  H��$�	  H��$�	  H��$`  H�$�    H��$�  H�\$H��$�  H�\$H��$   H�\$H��$  H��$�  H��H�� ��  H�� ��  H��$�	  W��    G�H��$�	  H��H�-    H�+H��$`  H�kH��$x  H�kH�KH��$h  H�k H��$p  H�k(H��$  H�k0H��$�  H�k8H��$�	  H�k@H��$`  H�� �Z  H�^ H�H�$H�KH�L$�D$H��$�  H����\$�� t郣��H��$�  H��$   H��$  H��$h  1�H��$`  H��$`  H��$X  H��$`  H9���   H��H��$�  H�� ��  H�	H�kH��$  H��$P  H��$X  H��$�  H�$H��$�  H�l$�D$ H��$�  H����\$�� t�ʢ��H��$�  H��$  H��H��H��$`  H9��j���H��$`  H�[(H�� ��  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hH�-    H�h H�-    H�h(HǄ$8     HǄ$@     H��$`  H�� ��  H�k H��$0  H�D$H�l$H�-    H�,$�    H��$0  H��$p  H�� H�kH��$h  �=     �:  H�+H��$`  H�$H��$0  H�\$H��$8  H�\$H��$@  H�\$�    H�L$ H�D$(H��$`  H�$H��$`  H�L$H��$h  H�D$�    �\$H�ـ� ��$�   ��  H��$�  H��H�� ��  H��$H  H�� �|  H�    H�$�    H�D$H�� �V  HǄ$`     HǄ$h     H��$`  H�� �%  H�k H��$X  H�D$H�l$H�-    H�,$�    H��$X  H��$H  H��H�kH��$@  �=     ��  H�+H��$`  H�$H��$X  H�\$H��$`  H�\$H��$h  H�\$�    H�L$ H�D$(H��$`  H�$H��$P  H�L$H��$X  H�D$�    ��$�   �\$H�؈�$�   �� ��  < ��  H��$`  H��$�	  H��$h  H��$�	  H��$�  H��$   H��$  H��$h  1�H��$`  H��$  H��$X  H��$  H9��Q  H��$�  H�� �
  H�H�hH��$`  H��$P  H��$�  H��$X  H��$�  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hH�-    H�h H�-    H�h(HǄ$x     HǄ$�     H��$p  H��$�  H�hH��$�  �=     �)  H�(H��$p  H��H�� H�kH��$h  �=     ��  H�+H��$`  H�$H�D$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$`  H�$H��$�  H�L$H��$�  H�D$�    �\$H�ـ� ��$�   �V  H��$�  H��H�� �@  H��$H  H�� �.  H�    H�$�    H�D$H�� �  HǄ$x     HǄ$�     H��$p  H��$�  H�hH��$�  �=     ��  H�(H��$H  H��H��H�kH��$@  �=     �f  H�+H��$`  H�$H�D$H��$x  H�\$H��$�  H�\$�    H�L$ H�D$(H��$`  H�$H��$P  H�L$H��$X  H�D$�    ��$�   �\$��$�   �� �d  ��$�    �V  H��$�	  H��$�	  H��$�	  H��H��H9���  H��$�	  H��H��Hk�H�H��$�  H�kH��$�  �=     ��  H�+H��$�  H��$`  H��H��H��$  H9������1�H��$�  H��$�  H��$�  H�    H��$�  HǄ$�     H��$�	  H��$�	  H��$�	  H��$h  1�H��$`  H��$  H��$X  H��$  H9���  H��$�  H�� ��
  H�H�hH��$`  H��$P  H��$X  H��$P  H��$�  H��$X  H��$�  1�H��$p  H��$x  H��$p  H�� �b
  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     ��	  H�CH��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�\$(H��$P  H�\$0H��$X  H��$�  H��$�  H��$�  H��H��H9���  H��$�  H��H��Hk�H�H��$X  H�kH��$P  �=     ��  H�+H�    H��$�  HǄ$�     H��$�  H��$`  H��H��H��$  H9�����H��$�	  H�� ��  1�H��$@  H��$H  H��$@  H�� ��  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�	  H�\$H�D$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     ��  H�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�\$(H��$P  H�\$0H��$X  H��$�  H��$�  H��$�  H��H��H9��  H��$�  H��H��Hk�H�H��$X  H�kH��$P  �=     ��  H�+H�    H��$�  HǄ$�     H��$�	  H��$�	  H��$�	  H��$�  1�H��$x  H��$`  H��$p  H��$`  H9���  H��H��$�  H�� �G  H�	H�kH��$  H��$P  H��$X  H��$p  H��$�  H��$x  H��$�  1�H��$0  H��$8  H��$0  H�� ��  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     �N  H�CH��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�\$(H��$P  H�\$0H��$X  H��$�  H��$�  H��$�  H��H��H9��n  H��$�  H��H��Hk�H�H��$X  H�kH��$P  �=     �%  H�+H�    H��$�  HǄ$�     H��$�  H��$  H��H��H��$`  H9��
���H��$�	  H�� uNH��$�  H��$�  H��$�  H��H��H9��T  H��$�  H��H��Hk�H�H�-    H�+H�C   H��$h  H��$�  H��$p  H��$�  H��$�  H�$H��$�  H�\$H��$�  H�\$H�    H�\$H�D$    �    H�\$(H��$�  H�\$0H��$�  1�H��$�  H��$�  H��$�  H��$�  H��$�  H�� �x  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     ��   H�CH�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$`  H�H��$h  �=     uvH�CH�    H�$H�D$$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$  H��$�  H��$�  H��$�  H��X  �L�CL�$H�D$�    �w���L�CL�$H�D$�    ���������H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  �^���H�$H�l$�    �����H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  �D���L�CL�$H�D$�    ��������������H�$H�l$�    �$���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  ����L�CL�$H�D$�    �������t���H��$�  H��$�  H��$�  H��H��H9�w,H��$�  H��H��Hk�H�H�-    H�+H�C   �a���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  �H�$H�l$�    �F���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  ����L�CL�$H�D$�    ���������� �-���H�$H�l$�    �`���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�	  H��$�	  H��$�	  �����H��$  H��$�  H�kH��$�  �=     uHH�+H��$  H��$�  H�kXH��$�  �=     u	H�kP�����L�CPL�$H�l$�    �ޏ��H�$H�l$�    �H�$H�l$�    H��$p  ����H�$H�l$�    H��$p  �<���� �����Ƅ$�    �����H�$H�l$�    H��$p  ����H�$H�l$�    H��$p  ����� �����H��$  H��$h  H�kH��$`  �=     udH�+H��$  H��   @���   H��$`  H�� t9H�k H��$  H�� t#L�CPL�D$H�l$H�-    H�,$�    �Ǝ����ى��H�$H�l$�    �H�$H�l$�    �1���������� ����1���$�   ����H�$H�l$�    ������Y�����;��������1������    1�����1�銉���    1��|���H��   �p���1������    1��ڈ��H��   �Έ��1��6���H��   �*���1��և����j���H��$X  H����   H�$H�D$H�-    H�l$H�D$   �    H��$`  �\$ �� ��   H�$    H�    H�\$H�D$
   H�� tmH�XH�|$H�H�H�KH�OH�    H�\$(H�D$0   H�|$8H�H�H�HH�OH��$P  H�\$HH��$X  H�\$P�    H�T$XH�L$`������ �H��$h  H��$�  H��$p  H��$�  1�H��$�  H��$�  H��$�  H��$�  H��$�  H�� ��  HǄ$�     HǄ$�     H��$�  H�    H�$H��$�  H�\$H�D$    �    H�L$H�D$ H��$�  H��$`  H�H��$h  �=     �  H�CH�    H�$H��$`  H�\$H�|$ ��   H�D$HH�D$    �    H�L$H�D$ H��$�  H��H��$`  H�H��$h  �=     usH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H��$   H��$(  H�\$(H��$0  H�\$0H��$8  �F���L�CL�$H�D$�    �z����%    �$���L�CL�$H�D$�    �������f���������鲂��L�@@L�$H�l$�    H��$�  靀����]����    �����

      \�  runtime.duffzero   ~�  runtime.duffzero   �  type."".Package   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  Tgo.string."import %q: invalid import path"   �  fmt.Errorf   �  .runtime.writebarrierptr   �
  go.string."_"   �  *runtime.concatstring2   �  go.string."gc"   �   runtime.eqstring   �   go.string."pkg/"   �  go.string."_"   �  *runtime.concatstring5   �  4"".(*Context).Import.func1   �       �  go.string."."   �   runtime.eqstring   �  go.string.".."   �   runtime.eqstring   �  go.string."./"   �   runtime.eqstring   �  go.string."../"   �   runtime.eqstring   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  vgo.string."import %q: import relative to unknown directory"   �  fmt.Errorf   �  .runtime.writebarrierptr   �   ."".(*Context).isAbsPath   �   type.[2]string   �   "runtime.newobject   �! (runtime.writeBarrier   �" (runtime.writeBarrier   �#  ,"".(*Context).joinPath   �$ (runtime.writeBarrier   �$  :"".(*Context).Import.func2·f   �$  type.[2]string   �%  "runtime.newobject   �%  """.statictmp_0250   �% """.statictmp_0250   �%  """.statictmp_0250   �%0 """.statictmp_0250   �&  type.string   �'  (runtime.typedmemmove   �'  ,"".(*Context).joinPath   �)  ."".(*Context).hasSubdir   �*       �+ (runtime.writeBarrier   �,  type.string   �,  (runtime.typedmemmove   �,  type.[2]string   �,  "runtime.newobject   �-  """.statictmp_0325   �- """.statictmp_0325   �-  """.statictmp_0325   �-0 """.statictmp_0325   �.  type.string   �.  (runtime.typedmemmove   �/  ,"".(*Context).joinPath   �0 (runtime.writeBarrier   �0  type.[2]string   �0  "runtime.newobject   �1  """.statictmp_0328   �1 """.statictmp_0328   �1  """.statictmp_0328   �10 """.statictmp_0328   �2  type.string   �2  (runtime.typedmemmove   �3  ,"".(*Context).joinPath   �4 (runtime.writeBarrier   �4  type.[2]string   �5  "runtime.newobject   �5  """.statictmp_0331   �5 """.statictmp_0331   �5  """.statictmp_0331   �50 """.statictmp_0331   �6  type.string   �7  (runtime.typedmemmove   �8  ,"".(*Context).joinPath   �8 (runtime.writeBarrier   �9  type.[2]string   �9  "runtime.newobject   �:  type.string   �;  (runtime.typedmemmove   �; (runtime.writeBarrier   �<  ,"".(*Context).joinPath   �= (runtime.writeBarrier   �=  type.[2]string   �>  "runtime.newobject   �?  type.string   �?  (runtime.typedmemmove   �@ (runtime.writeBarrier   �A  ,"".(*Context).joinPath   �B (runtime.writeBarrier   �E  *"".(*Context).readDir   �H  Ftype.map[string][]go/token.Position   �I  runtime.makemap   �I  Ftype.map[string][]go/token.Position   �J  runtime.makemap   �J  Ftype.map[string][]go/token.Position   �K  runtime.makemap   �L�  runtime.duffzero   �L  (type.map[string]bool   �M  runtime.makemap   �N  *type.go/token.FileSet   �N  "runtime.newobject   �N�  runtime.duffzero   �S       �W  "type."".NoGoError   �W  "runtime.newobject   �X  type.string   �X  (runtime.typedmemmove   �X  6go.itab.*"".NoGoError.error   �Z  $type.*"".NoGoError   �Z  type.error   �Z  6go.itab.*"".NoGoError.error   �Z   runtime.typ2Itab   �[�  runtime.duffzero   �[  (type.map[string]bool   �\  &runtime.mapiterinit   �^ (runtime.writeBarrier   �_  &runtime.mapiternext   �`  sort.Strings   �`  "".cleanImports   �a (runtime.writeBarrier   �b (runtime.writeBarrier   �c  "".cleanImports   �d (runtime.writeBarrier   �e (runtime.writeBarrier   �e  "".cleanImports   �g (runtime.writeBarrier   �g (runtime.writeBarrier   �i  type.[]string   �j  &runtime.growslice_n   �k  type.string   �m  ,runtime.typedslicecopy   �n (runtime.writeBarrier   �o  sort.Strings   �p  .runtime.writebarrierptr   �p  $runtime.panicslice   �p  $runtime.panicslice   �q  .runtime.writebarrierptr   �q  .runtime.writebarrierptr   �r  .runtime.writebarrierptr   �s  .runtime.writebarrierptr   �s  .runtime.writebarrierptr   �t  .runtime.writebarrierptr   �t  .runtime.writebarrierptr   �t  type.[]string   �u  "runtime.growslice   �v (runtime.writeBarrier   �v  .runtime.writebarrierptr   �w       �x  "".nameExt   �z  4"".(*Context).Import.func4   �|  ."".(*Context).matchFile   �       ��  go.string.".go"   ؀   runtime.eqstring   �� (runtime.writeBarrier   ҂  .runtime.writebarrierptr   �  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  go.string.".hh"   ҆  "runtime.cmpstring   ��  go.string.".h"   ��  "runtime.cmpstring   ��  go.string.".S"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ؋  type.[]string   ��  "runtime.growslice   ��  go.string.".c"   ��   runtime.eqstring   ȏ (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ̐  "runtime.growslice   ڑ (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  go.string.".h"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   Е  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]uint8   ��  runtime.convT2E   ֚  &go/parser.ParseFile   ��       ֝  2go.string."documentation"   ��   runtime.eqstring   ğ (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   Ƞ  "runtime.growslice   ֡ (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  (go.string."_test.go"   �   runtime.eqstring   ��  "go.string."_test"   ��   runtime.eqstring   �� (runtime.writeBarrier   ܯ  6go/ast.(*CommentGroup).Text   ̰  go/doc.Synopsis   ı (runtime.writeBarrier   ܲ  ("".findImportComment   ��  strconv.Unquote   ��  type.string   �  runtime.convT2E   �� (runtime.writeBarrier   �  type.int   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  \go.string."%s:%d: cannot parse import comment"   ��  fmt.Errorf   ��       ڿ  (type.*go/ast.GenDecl   ��  go.string."cgo"   ��  (type.map[string]bool   ��  $runtime.mapassign1   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  .type.*go/ast.ImportSpec   ��  strconv.Unquote   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  vgo.string."%s: parser returned invalid quoted string: <%s>"   ��  log.Panicf   ��  Ftype.map[string][]go/token.Position   ��  4runtime.mapaccess1_faststr   ��  8go/token.(*FileSet).Position   �� (runtime.writeBarrier   ��  Ftype.map[string][]go/token.Position   ��  $runtime.mapassign1   ��  go.string."C"   ��   runtime.eqstring   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  ^go.string."use of cgo in test %s not supported"   ��  fmt.Errorf   ��       ��  .runtime.writebarrierptr   ��  *"".(*Context).saveCgo   ��       ��  .runtime.writebarrierptr   ��  0type.[]go/token.Position   ��  "runtime.growslice   ��  Ftype.map[string][]go/token.Position   ��  4runtime.mapaccess1_faststr   Ȅ  8go/token.(*FileSet).Position   � (runtime.writeBarrier   ��  Ftype.map[string][]go/token.Position   �  $runtime.mapassign1   ��  .runtime.writebarrierptr   ��  0type.[]go/token.Position   ։  "runtime.growslice   ʌ  Ftype.map[string][]go/token.Position   ��  4runtime.mapaccess1_faststr   ֐  8go/token.(*FileSet).Position   �� (runtime.writeBarrier   ��  Ftype.map[string][]go/token.Position   �  $runtime.mapassign1   ��  .runtime.writebarrierptr   ��  0type.[]go/token.Position   �  "runtime.growslice   �  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��   runtime.eqstring   ���  runtime.duffzero   ��  type.string   ��  runtime.convT2E   � (runtime.writeBarrier   ��  type.string   ģ  runtime.convT2E   �� (runtime.writeBarrier   Ƥ  type.string   ��  runtime.convT2E   � (runtime.writeBarrier   ��  type.string   Ħ  runtime.convT2E   �� (runtime.writeBarrier   Ƨ  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  vgo.string."found import comments %q (%s) and %q (%s) in %s"   ��  fmt.Errorf   �       ��  .runtime.writebarrierptr   ܫ  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �  .runtime.writebarrierptr   ȭ  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �   runtime.eqstring   ��  8type."".MultiplePackageError   ��  "runtime.newobject   ��  type.string   ��  (runtime.typedmemmove   α  type.[2]string   �  "runtime.newobject   ��  type.string   ��  (runtime.typedmemmove   � (runtime.writeBarrier   ڴ (runtime.writeBarrier   ��  type.[2]string   ��  "runtime.newobject   �� (runtime.writeBarrier   �� (runtime.writeBarrier   ط (runtime.writeBarrier   ��  Lgo.itab.*"".MultiplePackageError.error   ¹       � (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   �  "runtime.growslice   �� (runtime.writeBarrier   Ľ  .runtime.writebarrierptr   ��  :type.*"".MultiplePackageError   ��  type.error   ��  Lgo.itab.*"".MultiplePackageError.error   ƾ   runtime.typ2Itab   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  $runtime.panicslice   ��  $runtime.panicslice   ��  $runtime.panicslice   ��  go.string.".s"   ��  "runtime.cmpstring   ��  go.string.".m"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  go.string.".s"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  go.string.".cc"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  go.string.".hh"   ��   runtime.eqstring   ��   go.string.".hpp"   ��  "runtime.cmpstring   ��   go.string.".cpp"   ��   runtime.eqstring   ��   go.string.".cxx"   ��   runtime.eqstring   ��   go.string.".hpp"   ��   runtime.eqstring   ��  "go.string.".swig"   ��  "runtime.cmpstring   ��   go.string.".hxx"   ��   runtime.eqstring   ��  "go.string.".swig"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  "go.string.".syso"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  (go.string.".swigcxx"   ��   runtime.eqstring   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  ("".(*Context).gopath   ��  type.[2]string   ��  "runtime.newobject   ��  """.statictmp_0257   �� """.statictmp_0257   ��  """.statictmp_0257   ��0 """.statictmp_0257   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  ."".(*Context).hasSubdir   ��       ��  type.[3]string   ��  "runtime.newobject   ��  """.statictmp_0260   �� """.statictmp_0260   ��  """.statictmp_0260   ��0 """.statictmp_0260   ��@ """.statictmp_0260   ��P """.statictmp_0260   ��  type.string   ��  (runtime.typedmemmove   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  &"".(*Context).isDir   �� (runtime.writeBarrier   ҁ  .runtime.writebarrierptr   Ą  type.[3]string   ք  "runtime.newobject   �  """.statictmp_0267   �� """.statictmp_0267   ��  """.statictmp_0267   ��0 """.statictmp_0267   ą@ """.statictmp_0267   څP """.statictmp_0267   ֆ (runtime.writeBarrier   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  &"".(*Context).isDir   � (runtime.writeBarrier   ��  .runtime.writebarrierptr   ΋ (runtime.writeBarrier   �� (runtime.writeBarrier   ܌  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  $runtime.panicslice   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ڐ  .runtime.writebarrierptr   ʑ  go.string."/"   ��   runtime.eqstring   ��  type.string     runtime.convT2E   �� (runtime.writeBarrier   ��  dgo.string."import %q: cannot import absolute path"   ��  fmt.Errorf   ��  .runtime.writebarrierptr   �  ("".(*Context).gopath   ���  runtime.duffzero   ֛  4"".(*Context).Import.func3   ��       �       ��  type.[3]string   ��  "runtime.newobject   ��  """.statictmp_0282   Ԣ """.statictmp_0282   �  """.statictmp_0282   ��0 """.statictmp_0282   ��@ """.statictmp_0282   ��P """.statictmp_0282   ¤  type.string   Ԥ  (runtime.typedmemmove   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  &"".(*Context).isDir   ��  type.[2]string   ��  "runtime.newobject   ک  type.string   �  (runtime.typedmemmove   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  ("".(*Context).isFile   ܯ  type.[3]string   �  "runtime.newobject   ��  """.statictmp_0291   �� """.statictmp_0291   ��  """.statictmp_0291   ư0 """.statictmp_0291   ܰ@ """.statictmp_0291   �P """.statictmp_0291   � (runtime.writeBarrier   Ĳ (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  &"".(*Context).isDir   ��  type.[2]string   µ  "runtime.newobject   Զ (runtime.writeBarrier   �� (runtime.writeBarrier   ��  ,"".(*Context).joinPath   ��  ("".(*Context).isFile   �� (runtime.writeBarrier   ��  <go.string."\t%s (vendor tree)"   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  fmt.Sprintf   �� (runtime.writeBarrier   ��   go.string."\t%s"   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  >go.string."\t%s (from $GOROOT)"   ��  fmt.Sprintf   �� (runtime.writeBarrier   ��  >go.string."\t%s (from $GOPATH)"   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  fmt.Sprintf   �� (runtime.writeBarrier   ��   go.string."\t%s"   ��  >go.string."\t($GOPATH not set)"   ��  go.string."\n"   ��  strings.Join   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  bgo.string."cannot find package %q in any of:\n%s"   ��  fmt.Errorf   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   ��  .runtime.writebarrierptr   ��  >go.string."\t($GOROOT not set)"   ��  type.[]string   ��  "runtime.growslice   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  type.[]string   ��  "runtime.growslice   �� (runtime.writeBarrier   �� (runtime.writeBarrier   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �� (runtime.writeBarrier   ��  type.string   ��  (runtime.typedmemmove   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  $runtime.panicslice   ��  $runtime.panicslice   ��  $runtime.panicslice   ��  "go.string."gccgo"   ��   runtime.eqstring   ��  ,go.string."pkg/gccgo_"   ��  go.string."_"   ��  *runtime.concatstring5   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  type.string   ��  runtime.convT2E   �� (runtime.writeBarrier   ��  Tgo.string."import %q: unknown compiler %q"   ��  fmt.Errorf   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   ��  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   ��-  �"".autotmp_0408  type.int "".autotmp_0407  type.[]string "".autotmp_0406  type.[]string "".autotmp_0405  Ftype.map[string][]go/token.Position "".autotmp_0404  type.[]string "".autotmp_0403  Ftype.map[string][]go/token.Position "".autotmp_0402  type.[]string "".autotmp_0401 �$Ftype.map[string][]go/token.Position "".autotmp_0400  type.[]string "".autotmp_0399  type.*uint8 "".autotmp_0398 �$$type.*"".NoGoError "".autotmp_0397  "type.interface {} "".autotmp_0396  (type.[1]interface {} "".autotmp_0394  *type.*[1]interface {} "".autotmp_0393  &type.[]interface {} "".autotmp_0392  "type.go/token.Pos "".autotmp_0391  "type.go/token.Pos "".autotmp_0390  "type.go/token.Pos "".autotmp_0389  "type.go/token.Pos "".autotmp_0388  "type.go/token.Pos "".autotmp_0387 �)"type.go/token.Pos "".autotmp_0386  "type.interface {} "".autotmp_0385  "type.interface {} "".autotmp_0384 �(type.[2]interface {} "".autotmp_0382  *type.*[2]interface {} "".autotmp_0381  &type.[]interface {} "".autotmp_0380 � type.go/ast.Spec "".autotmp_0379 �#"type.*go/ast.Spec "".autotmp_0378 �)type.int "".autotmp_0377 �)type.int "".autotmp_0376 � type.go/ast.Decl "".autotmp_0375 �#"type.*go/ast.Decl "".autotmp_0374  type.int "".autotmp_0373  type.int "".autotmp_0372  "type.interface {} "".autotmp_0371  "type.interface {} "".autotmp_0370  "type.interface {} "".autotmp_0369  "type.interface {} "".autotmp_0368  "type.interface {} "".autotmp_0367 �(type.[5]interface {} "".autotmp_0365 �#*type.*[5]interface {} "".autotmp_0364  &type.[]interface {} "".autotmp_0363  type.string "".autotmp_0362  "type.interface {} "".autotmp_0361  "type.interface {} "".autotmp_0360  (type.[2]interface {} "".autotmp_0358  *type.*[2]interface {} "".autotmp_0357  &type.[]interface {} "".autotmp_0356 �#type.*uint8 "".autotmp_0355  type.*[2]string "".autotmp_0354  type.[]string "".autotmp_0353  type.*[2]string "".autotmp_0352  type.[]string "".autotmp_0351 �#:type.*"".MultiplePackageError "".autotmp_0350 �type.string "".autotmp_0349  type.bool "".autotmp_0348  type.bool "".autotmp_0347  type.string "".autotmp_0346 �	�type.struct { F uintptr; badGoError *error; p *"".Package; name string } "".autotmp_0345 �#�type.*struct { F uintptr; badGoError *error; p *"".Package; name string } "".autotmp_0344 � type.os.FileInfo "".autotmp_0343 �#"type.*os.FileInfo "".autotmp_0342  type.int "".autotmp_0341  type.int "".autotmp_0340 �#,type.*go/token.FileSet "".autotmp_0339  ,type.*go/token.FileSet "".autotmp_0338 �6type.map.bucket[string]bool "".autotmp_0337 �0type.map.hdr[string]bool "".autotmp_0336  type.*[2]string "".autotmp_0335  type.[]string "".autotmp_0334  type.*[2]string "".autotmp_0333  type.[]string "".autotmp_0332  type.*[2]string "".autotmp_0330  type.[]string "".autotmp_0329  type.*[2]string "".autotmp_0327  type.[]string "".autotmp_0326  type.*[2]string "".autotmp_0324  type.[]string "".autotmp_0323  "type.interface {} "".autotmp_0322  "type.interface {} "".autotmp_0321 �
(type.[2]interface {} "".autotmp_0319  *type.*[2]interface {} "".autotmp_0318  &type.[]interface {} "".autotmp_0317  "type.interface {} "".autotmp_0316 �(type.[1]interface {} "".autotmp_0314  *type.*[1]interface {} "".autotmp_0313  &type.[]interface {} "".autotmp_0312  type.string "".autotmp_0311  type.*string "".autotmp_0310  type.int "".autotmp_0309  type.int "".autotmp_0308  "type.interface {} "".autotmp_0307 �(type.[1]interface {} "".autotmp_0305  *type.*[1]interface {} "".autotmp_0304  &type.[]interface {} "".autotmp_0303  "type.interface {} "".autotmp_0302  (type.[1]interface {} "".autotmp_0300  *type.*[1]interface {} "".autotmp_0299  &type.[]interface {} "".autotmp_0298  type.string "".autotmp_0297  type.*string "".autotmp_0296  type.int "".autotmp_0295  type.int "".autotmp_0294  type.*[2]string "".autotmp_0293  type.[]string "".autotmp_0292  type.*[3]string "".autotmp_0290  type.[]string "".autotmp_0289  type.string "".autotmp_0288  type.*string "".autotmp_0287  type.int "".autotmp_0286  type.int "".autotmp_0285  type.*[2]string "".autotmp_0284  type.[]string "".autotmp_0283  type.*[3]string "".autotmp_0281  type.[]string "".autotmp_0280  type.string "".autotmp_0279  type.*string "".autotmp_0278  type.int "".autotmp_0277  type.int "".autotmp_0276 ��type.struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } } "".autotmp_0274  "type.interface {} "".autotmp_0273  (type.[1]interface {} "".autotmp_0271  *type.*[1]interface {} "".autotmp_0270  &type.[]interface {} "".autotmp_0269  type.bool "".autotmp_0268  type.*[3]string "".autotmp_0266 �type.[]string "".autotmp_0265  type.string "".autotmp_0264 �"type.*string "".autotmp_0263 �)type.int "".autotmp_0262  type.int "".autotmp_0259  type.[]string "".autotmp_0258  type.*[2]string "".autotmp_0256 �type.[]string "".autotmp_0255  type.string "".autotmp_0254 �"type.*string "".autotmp_0253  type.int "".autotmp_0252  type.int "".autotmp_0251  type.*[2]string "".autotmp_0249  type.[]string "".autotmp_0247 �type.[]string "".autotmp_0246  "type.interface {} "".autotmp_0245  (type.[1]interface {} "".autotmp_0243  *type.*[1]interface {} "".autotmp_0242  &type.[]interface {} "".autotmp_0241  type.bool "".autotmp_0240  type.bool "".autotmp_0239  type.bool "".autotmp_0238 ��type.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } "".autotmp_0236  "type.interface {} "".autotmp_0235  "type.interface {} "".autotmp_0234 �
(type.[2]interface {} "".autotmp_0231  &type.[]interface {} "".autotmp_0230 �type.string "".autotmp_0229 �'type.[32]uint8 "".autotmp_0228 �"type.interface {} "".autotmp_0227 �(type.[1]interface {} "".autotmp_0224 �&type.[]interface {} "".autotmp_0223 �" type.*"".Package "".autotmp_0222  type.int "".autotmp_0221 �2type.map.iter[string]bool "".autotmp_0220 �"(type.map[string]bool "".autotmp_0219  $type.*"".NoGoError "".autotmp_0218  type.int "".autotmp_0217  type.int "".autotmp_0216  type.int "".autotmp_0215  type.int "".autotmp_0214 �+type.bool "".autotmp_0213  type.string "".autotmp_0212 �)type.int "".autotmp_0211  type.error "".autotmp_0210  type.string "".autotmp_0209  0type.[]go/token.Position "".autotmp_0208  ,type.go/token.Position "".autotmp_0207  0type.[]go/token.Position "".autotmp_0206  type.string "".autotmp_0205  type.string "".autotmp_0204  0type.[]go/token.Position "".autotmp_0203  ,type.go/token.Position "".autotmp_0202  0type.[]go/token.Position "".autotmp_0201  type.string "".autotmp_0200  type.string "".autotmp_0199 �0type.[]go/token.Position "".autotmp_0198 �	,type.go/token.Position "".autotmp_0197 �0type.[]go/token.Position "".autotmp_0196  type.string "".autotmp_0195  type.string "".autotmp_0194  type.string "".autotmp_0193  type.string "".autotmp_0192 �".type.*go/ast.ImportSpec "".autotmp_0191 �$type.[]go/ast.Spec "".autotmp_0190 �"(type.*go/ast.GenDecl "".autotmp_0189 �$type.[]go/ast.Decl "".autotmp_0188  type.error "".autotmp_0187 �type.string "".autotmp_0186  type.string "".autotmp_0185  type.string "".autotmp_0184  type.error "".autotmp_0183 �(type.int "".autotmp_0182  type.string "".autotmp_0181 �type.string "".autotmp_0180  type.string "".autotmp_0179  :type.*"".MultiplePackageError "".autotmp_0178  type.int "".autotmp_0177  type.int "".autotmp_0176 �type.string "".autotmp_0175 �(type.int "".autotmp_0174 �(type.int "".autotmp_0173 �(type.int "".autotmp_0172  type.int "".autotmp_0171  type.int "".autotmp_0170  type.string "".autotmp_0169 �(type.int "".autotmp_0168 �(type.int "".autotmp_0167 �(type.int "".autotmp_0166  type.int "".autotmp_0165  type.int "".autotmp_0164 �type.[]uint8 "".autotmp_0163  type.bool "".autotmp_0162 �$type.[]os.FileInfo "".autotmp_0161  type.string "".autotmp_0160  type.string "".autotmp_0159  type.string "".autotmp_0158  type.string "".autotmp_0157  type.string "".autotmp_0156  type.error "".autotmp_0155 �type.string "".autotmp_0154  type.string "".autotmp_0153  type.int "".autotmp_0152  type.string "".autotmp_0151  type.string "".autotmp_0150  type.[]string "".autotmp_0149  type.string "".autotmp_0148  type.string "".autotmp_0147  type.string "".autotmp_0146  type.[]string "".autotmp_0145  type.bool "".autotmp_0144  type.string "".autotmp_0143  type.[]string "".autotmp_0142  type.bool "".autotmp_0141  type.string "".autotmp_0140  type.bool "".autotmp_0139  type.[]string "".autotmp_0138  type.bool "".autotmp_0137  type.error "".autotmp_0136  type.string "".autotmp_0135  type.string "".autotmp_0134  type.int "".autotmp_0133  type.int "".autotmp_0132  type.int "".autotmp_0131  type.bool "".autotmp_0130 �type.[]string "".autotmp_0129  type.[]string "".autotmp_0128  type.bool "".autotmp_0127  type.bool "".autotmp_0126  type.[]string "".autotmp_0125  type.bool "".autotmp_0124  type.string "".autotmp_0123  type.bool "".autotmp_0122  type.error "".autotmp_0121  type.string "".autotmp_0120  type.string "".autotmp_0119  type.int "".autotmp_0118  type.int "".autotmp_0117  type.int "".autotmp_0116  type.string "".autotmp_0115 �(type.int "".autotmp_0114 �'type.int "".autotmp_0113 �'type.int "".autotmp_0112  type.string "".autotmp_0111 �type.error "".autotmp_0110 �type.string "".~r0 �*"type.go/token.Pos go/ast.x·2 �&*type.*go/ast.BasicLit "".~r0 �*"type.go/token.Pos go/ast.x·2 �&$type.*go/ast.Ident "".~r0 �+"type.go/token.Pos go/ast.s·2 �%.type.*go/ast.ImportSpec "".~r0 �*"type.go/token.Pos go/ast.x·2 �&*type.*go/ast.BasicLit "".~r0 �+"type.go/token.Pos go/ast.x·2 �'$type.*go/ast.Ident "".~r0 �*"type.go/token.Pos go/ast.s·2 �&.type.*go/ast.ImportSpec "".~r0 �*"type.go/token.Pos go/ast.x·2 �&*type.*go/ast.BasicLit "".~r0 �*"type.go/token.Pos go/ast.x·2 �&$type.*go/ast.Ident "".~r0 �*"type.go/token.Pos go/ast.s·2 �%.type.*go/ast.ImportSpec "".~r0 �+type.bool "strings.suffix·3 � type.string strings.s·2 �!type.string "".~r0 �+type.bool "strings.suffix·3 � type.string strings.s·2 �!type.string "".~r0 �',type.*go/token.FileSet "strings.prefix·3 �type.string strings.s·2 �!type.string "strings.prefix·3 �type.string strings.s·2 �!type.string "strings.prefix·3 �type.string strings.s·2 � type.string "".path �type.string "".tag �"type.string "".err �type.error 
"".cg �$2type.*go/ast.CommentGroup "".err �type.error "".path �type.string "".quoted �type.string 
"".ok �+type.bool "".spec �%.type.*go/ast.ImportSpec "".dspec � type.go/ast.Spec 
"".ok �+type.bool "".d �$(type.*go/ast.GenDecl "".decl � type.go/ast.Decl "".isCgo �+type.bool "".err �type.error "".com �type.string "".line �*type.int "".qcom �type.string "".isXTest �+type.bool "".isTest �+type.bool "".pkg �type.string 
"".pf �%"type.*go/ast.File "".err �type.error "".filename �type.string "".data �type.[]uint8 "".match �+type.bool "".badFile �$ type.func(error) "".ext �type.string "".name �type.string "".d � type.os.FileInfo "".fset �$,type.*go/token.FileSet "".allTags �"(type.map[string]bool  "".xTestImported �&Ftype.map[string][]go/token.Position "".testImported �&Ftype.map[string][]go/token.Position "".imported �$Ftype.map[string][]go/token.Position &"".firstCommentFile �type.string "".firstFile �type.string "".Sfiles �type.[]string "".badGoError �type.error "".err �type.error "".dirs �$type.[]os.FileInfo "".dir �type.string "".dir �type.string "".format �type.string "".paths �type.[]string "".isDir �+type.bool "".dir �type.string "".root �type.string "".isDir �+type.bool "".dir �type.string "".root �type.string "".searchVendor �%8type.func(string, bool) bool "".gopath �type.[]string "".tried �~type.struct { vendor []string; goroot string; gopath []string } "".dir �type.string "".earlyRoot �type.string "".dir �type.string "".sub �type.string "".rootsrc �type.string "".root �type.string "".i �)type.int "".all �type.[]string "".sub �type.string "".root �type.string "".inTestdata �%,type.func(string) bool "".binaryOnly �+type.bool "".setPkga �%type.func() "".suffix � type.string "".pkgerr �type.error "".pkga �type.string  "".pkgtargetroot �type.string "".p �% type.*"".Package "".~r4 ptype.error "".~r3 ` type.*"".Package "".mode P$type."".ImportMode "".srcDir 0type.string "".path type.string "".ctxt   type.*"".Context �"�-��-�-��-�-��-�-S�-�-��-�-��-�-��-�-��-�-���-�-�#�-�-��-
 
�� ��q[�l"[�
���9���%>������88m8$888���(0�8r��d$7���
!�;0
	0((��4@��&!(S\+,+,�� SXYZYZVS\;<;<�C\MNMN�,�&}�.S\�������%- -�RR��T@PZ\�����\�����\�����\�����\�����]�T,
.R��S�%&1m&;�����55) ����>��6\�5T!MZS\GHGH�
C\STST�S\ABAB�
C.AZ�C.AZOC\_`_`�
S\qrqr�C\efef�e-((� ����/������/����())����6	DT��B@ �6Bvo5no(�3� ��3�
`(|�(��(N�Vt	tJStV()<;<=J6(>RQ/Qg\!K�
�A
 �	 |�rD�q��R��rD7��8���8�8�8�h:�h�88�)��JK�������[QJ))!!!!	)k=O5��U})kl�)g�)kN}	)ko�u})k�
����� �E)k�)k�)k�)k�)k�*�����E�rG�i)���9���9���y��G�	|ioy��A7A.o	�)kN}	)kN�)kNN�N�}	)kN�)kN}	)k<((9���1�h5S��5S�46)��rD_�*�Z�h5�h����{�v�{�����DG@	)D!)D=	)D!y)�38J�-+*/&+�	���AO# Tgclocals·3b32eac464325adfcb2e0feeafb27ba3 Tgclocals·5391224ff1aeba9fa698864a89676656   :$GOROOT/src/go/build/build.go�"".hasGoFiles  �  �dH�%    H�D$�H;A��  H���   H��$�   H�$H��$�   H�\$H��$�   H�\$�    H�T$H�D$ H�L$(H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$@H��$�   H��H�l$@H9��&  H�D$PH�� �6  H�H�hH�L$HH��$�   H��$�   H��$�   H�,$H�T$xH�Z ���\$�� ��   H��$�   H�$H�\$xH�[8��H�|$H�L$H�|$XH�5    H�t$hH��   H�L$`H�D$pH9���   H��H)�H��H9���   H)�I��H�� tM�H9�usL��$�   L�$H��$�   H�l$H�t$H�D$�    �\$ H��< tƄ$�   H���   �H�D$PH�L$HH��H��H�l$@H9������Ƅ$�    H���   �1���    1�뮉 ������    �	������������
      �  *"".(*Context).readDir   �       �       �  go.string.".go"   �   runtime.eqstring   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0508 � type.os.FileInfo "".autotmp_0507 �"type.*os.FileInfo "".autotmp_0506 �type.int "".autotmp_0505 �type.int "".autotmp_0504  type.string "".autotmp_0498 type.string "".autotmp_0496 /$type.[]os.FileInfo "strings.suffix·3 �type.string strings.s·2 �type.string "".ent � type.os.FileInfo "".ents _$type.[]os.FileInfo "".~r2 0type.bool "".dir type.string "".ctxt   type.*"".Context ,����.��� � .�:s�
  E�%�% Tgclocals·14c16763214c88f6ebc22b4b638329b7 Tgclocals·80ce1eebd7f944e81966bdd86878cedc   :$GOROOT/src/go/build/build.go�("".findImportComment  �  �dH�%    H�D$�H;A��  H��   1�1�H��$�   H��$�   H��$�   H�$H��$�   H�\$H��$�   H�\$�    H�T$H�L$ H�D$(H�\$0H��$�   H�\$8H��$�   H�\$@H��$�   H�T$XH�$H�L$`H�L$H�D$hH�D$�    H�L$H�D$ H����  H�L$HH�$H�D$PH�D$H�-    H�l$H�D$   �    �\$ �� ��  H��$�   H�$H��$�   H�\$H��$�   H�\$�    H�L$0H�D$8H�T$@H�� ~GH�� �a  ��� �  H��H��H���  H��H��I��H�� tI��H��H��L��H�� �1�H�\$pH�\$xH��$�   H��$�   H�$H��$�   H�D$H��$�   H�T$H�    H�\$H�    H�\$ H�    H�\$(�    H��$�   H��$�   H��$�   �\$0�� ��  H�,$H�T$H�L$H�    H�\$H�    H�\$ H�    H�\$(�    H�D$0H�� }H��$�   H��$�   H��H9��Y  H���O  L��$�   H��H��H�� tI��H�\$xH��$�   L�D$pH�\$pH�$H�\$xH�\$H��$�   H�\$�    H�T$H�L$ H�D$(H�T$pH�$H�L$xH�L$H��$�   H�D$�    H�T$H�L$ H�D$(H�\$0H��$�   H�\$8H��$�   H�\$@H��$�   H�T$XH�$H�L$`H�L$H�D$hH�D$�    H�L$H�D$ H���8  H�L$HH�$H�D$PH�D$H�-    H�l$H�D$   �    H��$�   �\$ �� ��   H��$�   H��H)�H9���   L��$�   L��$�   L�$H��$�   H�\$H��$�   H�T$H�    H�\$H�    H�\$ H�    H�\$(�    H�\$0H��H��$�   H�$    H��$�   H�\$H��$�   H�\$H��$�   H�\$�    H�\$ H�H�$H�KH�L$�    H�L$H�D$H��$�   H��$�   H�ĸ   ��    1�H��$�   H��$�   HǄ$�       H�ĸ   ��    H�,$H�T$H�L$H�    H�\$H�    H�\$ H�    H�\$(�    �\$0�� �����H��$�   H��$�   H���8  L��$�   H��H��H�� tI��L��$�   L�$H��$�   H�\$H��$�   H�l$H�    H�\$H�    H�\$ H�    H�\$(�    H�D$0H�� }&1�H��$�   H��$�   HǄ$�       H�ĸ   �H��$�   H9���   L��$�   L�D$pL�$H�D$xH�D$H��$�   H�l$H�    H�\$H�    H�\$ H�    H�\$(�    �\$0�� t&1�H��$�   H��$�   HǄ$�       H�ĸ   ��F����    �    �    H�� v+���	u�����H�� v�������������    �    �    1�H��$�   H��$�   HǄ$�       H�ĸ   ��    �������������\
      �  "".parseWord   �  8runtime.slicebytetostringtmp   �  &go.string."package"   �   runtime.eqstring   �  "".parseWord   �  "".slashSlash   � "".slashSlash   �  "".slashSlash   �  bytes.HasPrefix   �  "".newline   � "".newline   �  "".newline   �	  bytes.Index   �  bytes.TrimSpace   �  "".parseWord   �  8runtime.slicebytetostringtmp   �  $go.string."import"   �   runtime.eqstring   �  "".newline   � "".newline   �  "".newline   �  bytes.Count   �  2runtime.slicebytetostring   �  "strings.TrimSpace   �  $runtime.panicslice   �  $runtime.panicslice   �  "".slashStar   � "".slashStar   �  "".slashStar   �  bytes.HasPrefix   �  "".starSlash   � "".starSlash   �  "".starSlash   �  bytes.Index   �  "".newline   � "".newline   �  "".newline   �  bytes.Contains   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `�  "".autotmp_0521  type.string "".autotmp_0520 �type.string "".autotmp_0519  type.string "".autotmp_0517 _type.[]uint8 "".autotmp_0514  type.int "".arg /type.[]uint8 "".comment �type.[]uint8 "".word �type.[]uint8 "".line Ptype.int "".s 0type.string "".data  type.[]uint8 H����,��������~� � ��3aq
:+u<J4[y~p&#E4T&S&?& 8 Y�]�����:� Tgclocals·adb3347b296419e60da36d67f8b7ce43 Tgclocals·423fcdc350b935457e47f75dd5e63926   :$GOROOT/src/go/build/build.go�*"".skipSpaceOrComment  �  �dH�%    H;a��  H��8H�t$PH�T$@H�L$H1�H�\$XH�\$`H�\$hH�� ~FH�� �s  �*@��
wV@��	uHH��H��H��r5H��H��I��H�� tI��H��H��L��H�� �H�T$XH�L$`H�t$hH��8��    @��
t���@��t�@�� t�@��/u�H�T$@H�$H�L$HH�L$H�t$PH�t$H�    H�\$H�    H�\$ H�    H�\$(�    H�l$HH�T$@H�L$P�\$0�� ��   H�$H�l$H�L$H�    H�\$H�    H�\$ H�    H�\$(�    H�D$0H�� }1�H�\$XH�\$`H�\$hH��8�H��H��H�l$HL�D$PH9�w9L�L$@H)�I)�I�� tM�H��L��L��H�� �����H�� ������    �    H�$H�l$H�L$H�    H�\$H�    H�\$ H�    H�\$(�    H�t$PH�T$@H�L$H�\$0�� ��   H��H��H����   H��H��I��H�� tI��L�D$@L�$H�\$HH�\$H�l$PH�l$H�    H�\$H�    H�\$ H�    H�\$(�    H�D$0H�� }1�H�\$XH�\$`H�\$hH��8�H�l$HL�D$PH��H��H9�w#L�L$@H)�I)�I�� tM�H��L��L���V����    �    �����    ������.
      �  $runtime.panicslice   �  "".slashSlash   � "".slashSlash   �  "".slashSlash   �  bytes.HasPrefix   �  "".newline   � "".newline   �  "".newline   �  bytes.Index   �  $runtime.panicindex   �  $runtime.panicslice   �  "".slashStar   � "".slashStar   �  "".slashStar   �  bytes.HasPrefix   �	  "".starSlash   �	 "".starSlash   �	  "".starSlash   �
  bytes.Index   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   `p  "".autotmp_0526  type.int "".autotmp_0525  type.bool "".~r1 0type.[]uint8 "".data  type.[]uint8 *pop�op�opLo � ��7'4-c<3
T%K4'(	  �� Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�"".parseWord  �  �dH�%    H;a�{  H��@1�1�1�H�\$xH��$�   H��$�   1�H�\$`H�\$hH�\$pH�\$HH�$H�\$PH�\$H�\$XH�\$�    H�T$H�L$ H�D$(H�T$HH�L$PH�D$XH�T$xH�$H��$�   H�L$H��$�   H�D$�    �D$H�\$ H�\$8�D$4�$�    H��$�   �L$4�\$�� u
��0|D��9?H�\$8L��$�   H��H9�w#L�L$xH)�I)�I�� tM�H��L��L���f����    ��_t�H�\$PH�l$XH)�H9�wLL�D$HH�l$pL�D$`H�\$hH�� u-1�H�\$`H�\$hH�\$p1�H�\$xH��$�   H��$�   H��@�H��@��    �    �h�����������
      �  *"".skipSpaceOrComment   �  .unicode/utf8.DecodeRune   �   unicode.IsLetter   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   ��  "".autotmp_0532  type.int "".size type.int "".r type.int32 "".rest `type.[]uint8 "".word 0type.[]uint8 "".data  type.[]uint8 &���� � @�C16,3!-	  `Fw� Tgclocals·b4015c155c4a804136b8d2d3fde81a78 Tgclocals·69c1753bd5f81501d95132d08af04464   :$GOROOT/src/go/build/build.go�."".(*Context).MatchFile  �  �dH�%    H;a��   H��x1�1�H��$�   H��$�   H��$�   H�$H��$�   H�\$H��$�   H�\$H��$�   H�\$H��$�   H�\$ �D$( H�D$0    �    �\$8��$�   H�\$hH��$�   H�\$pH��$�   H��x��    �M����������������
      �  ."".(*Context).matchFile   �  0runtime.morestack_noctxt   ��  
"".err `type.error "".match Ptype.bool "".name 0type.string "".dir type.string "".ctxt   type.*"".Context ��� � �+y 
 yG Tgclocals·a043b57aa077fd78befe739904a3c363 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�."".(*Context).matchFile  �<  �<dH�%    H��$8���H;A��  H��H  1�1�1�1�H��$�  H��$�  1�H��$�  H��$�  1�H��$�  H��$�  H��$�  Ƅ$�   L��$h  L�D$HH��$p  H�=    H��$�   H��   H�t$PH��$�   H9��K  H9��;  H9��+  L��$�   L�$H��$�   H�D$H�|$H�D$�    �\$ H��< ��  H��$h  H�|$hH��$p  H�5    H��$�   H��   H�L$pH��$�   H9���  H9���  H9���  H��$�   H�<$H��$�   H�D$H�t$H�D$�    �\$ H��< �K  H��$h  H�$H��$p  H�\$H�    H�\$H�D$   �    H��$h  H��$p  H�D$ H�� }H��H��H9���  H)�I��H�� tM� H��$�   L��$�   H��$P  H�$H�T$H�L$H��$�  H�\$�    �\$ �� uH��$P  �]A�� uH��H  �H��$�   H��$�   H��$�   H��|TH����  H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� �t  H��|TH����  H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� ��  H����  H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� ��  H�    H�$�    H�D$H�� �k  HǄ$     HǄ$      H��$  H��$`  H�hH��$X  �=     �  H�(H��$p  H��H��H�kH��$h  �=     ��  H�+H��$P  H�$H�D$H��$  H�\$H��$   H�\$�    H�L$ H�D$(H��$P  H�$H��$�  H�L$H��$�  H�D$�    L�T$L��$�   L�L$ L��$�   H�D$(H�\$0H��$�  H��$�  H�� tH��H  �H��$�  H�|$XH��$�  H�5    H�t$xH��   H�L$`H��$�   H9���  H��H)�H��H9���  H)�I��H�� tM�H9���  L��$�   L�$H��$�   H�l$H�t$H�D$�    L��$�   L��$�   �\$ H��< ��  H�    H�$L�T$L�L$�    H�\$H�H�$H�KH�L$�D$ H�D$    �    H�\$ H��$�  H�\$(H��$�  H�\$0H��$�  H�\$8H��$�  H�\$@H��$�  H��$�   H�$H��$�   H�[ ��H��$�  H�� ��  H��$�  H��$�   H��$�  H��$�   1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �]  HǄ$      HǄ$     H��$�   H�    H�$H��$�   H�\$H�D$    �    H�L$H�D$ H��$�   H��$�   H�H��$�   �=     ��   H�CH��$�  H�$H��$�  H�\$�    H�L$H�D$H��$�   H��H��$�   H�H��$�   �=     ufH�CH�    H�$H�D$   H��$�   H�\$H��$   H�\$H��$  H�\$ �    H�\$(H��$�  H�\$0H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H��$P  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    �\$(�� uH��$P  �]A�� uH��H  �Ƅ$�  H��H  �H�    H�$L�T$L�L$�    H�\$H�H�$H�KH�L$�    H�\$H��$�  H�\$H��$�  H�\$ H��$�  H�\$(H��$�  H�\$0H��$�  �*���1������    1�����H�$H�l$�    H��$  ����H�$H�l$�    H��$  ������ ����H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� � ���H��uAH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� �����H��H  �H��|TH����   H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� ��   H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� �(���H���E���H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� ����������H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� �����H�������H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� �>����`���H��|TH����  H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� ��  H��|TH����   H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� ��   H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� �6���H���S���H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� ���������H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� �����H�������H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� �L����n���H��|TH����   H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   H�\$ H�� ��   H��uIH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� �����H�������H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� �S����u���H��uUH��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� tƄ$�  H��H  �H������H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� �����������    H��H  �1������    1�����1�������    1�������    ���������̤
      �  go.string."_"   �   runtime.eqstring   �  go.string."."   �   runtime.eqstring   �  go.string."."   �  "strings.LastIndex   �  8"".(*Context).goodOSArchFile   �
  go.string.".go"   �
  "runtime.cmpstring   �  go.string.".h"   �  "runtime.cmpstring   �  go.string.".S"   �   runtime.eqstring   �  type.[2]string   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   �  ,"".(*Context).joinPath   �  ,"".(*Context).openFile   �  go.string.".go"   �   runtime.eqstring   �  type.io.Reader   �  runtime.convI2I   �  "".readImports   �       �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  runtime.convI2E   � (runtime.writeBarrier   �  .go.string."read %s: %v"   �  fmt.Errorf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  2"".(*Context).shouldBuild   �   type.io.Reader   �!  runtime.convI2I   �!  "".readComments   �"  $runtime.panicslice   �#  .runtime.writebarrierptr   �#  .runtime.writebarrierptr   �$  go.string.".c"   �$   runtime.eqstring   �%  go.string.".h"   �&   runtime.eqstring   �'  go.string.".s"   �'  "runtime.cmpstring   �(  go.string.".m"   �(   runtime.eqstring   �)  go.string.".s"   �)   runtime.eqstring   �*  go.string.".cc"   �+   runtime.eqstring   �,  go.string.".go"   �,   runtime.eqstring   �-   go.string.".hpp"   �-  "runtime.cmpstring   �.   go.string.".cpp"   �/  "runtime.cmpstring   �0  go.string.".hh"   �0   runtime.eqstring   �1   go.string.".cpp"   �1   runtime.eqstring   �2   go.string.".cxx"   �2   runtime.eqstring   �3   go.string.".hpp"   �4   runtime.eqstring   �5  "go.string.".swig"   �5  "runtime.cmpstring   �6   go.string.".hxx"   �6   runtime.eqstring   �7  "go.string.".swig"   �8   runtime.eqstring   �8  "go.string.".syso"   �9   runtime.eqstring   �:  (go.string.".swigcxx"   �:   runtime.eqstring   �;  $runtime.panicslice   �;  $runtime.panicslice   �;  $runtime.panicslice   �<  0runtime.morestack_noctxt   ��  J"".autotmp_0561  "type.interface {} "".autotmp_0560 �"type.interface {} "".autotmp_0559 ?(type.[2]interface {} "".autotmp_0556 �&type.[]interface {} "".autotmp_0555  type.bool "".autotmp_0553 otype.[]string "".autotmp_0552  type.string "".autotmp_0551  type.bool "".autotmp_0549  type.bool "".autotmp_0548 �type.string "".autotmp_0547  type.string "".autotmp_0544  type.int "".autotmp_0543  type.int "".autotmp_0542  type.int "".autotmp_0541  type.bool "".autotmp_0540  type.string "".autotmp_0539  type.int "".autotmp_0538  type.int "".autotmp_0537  type.int "".autotmp_0536 �type.string "strings.suffix·3 �type.string strings.s·2 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "".f �$type.io.ReadCloser "".ext �type.string "".err �type.error "".filename �type.string "".data �type.[]uint8 "".match ptype.bool "".allTags `(type.map[string]bool  "".returnImports Ptype.bool "".name 0type.string "".dir type.string "".ctxt   type.*"".Context ~"�������������������	��^��*� � ��n��H,C�S�W���2
`u	=�Z�����Z�K	K � ��~�����Tv4QMl
hOY�LSV�LSV�L_H Tgclocals·d644b00c61b0153799eb59e0efc3a880 Tgclocals·8464a0493338a790ce587fd837b5331f   :$GOROOT/src/go/build/build.go�"".cleanImports  �  �dH�%    H�D$�H;A�  H���   1�H��$�   H��$�   H��$�   H��$�   1�H9�tH�H��H�    H�$H�D$    H�D$�    H�\$H�\$PH�\$ H�\$XH�\$(H�\$`H��$�   H�|$hW�H����    H�    H�$H�D$H�\$hH�\$�    H�\$h1�H9���   H�\$hH�� �>  H�+H�l$@H�kH�l$HH�L$PH�D$XH�T$`H��H��H9���   H�\$XH��H��Hk�H�H�l$HH�kH�l$@�=     ��   H�+H�\$hH�$�    H�\$h1�H9��t���H�\$PH�$H�\$XH�\$H�\$`H�\$�    H�\$PH��$�   H�\$XH��$�   H�\$`H��$�   H��$�   H��$�   H���   �H�$H�l$�    �n���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�D$0H�T$8H��H��H�\$XH�T$`H�L$P�����������    �����
      �  type.[]string   �  "runtime.makeslice   ��  runtime.duffzero   �  Ftype.map[string][]go/token.Position   �  &runtime.mapiterinit   � (runtime.writeBarrier   �  &runtime.mapiternext   �  sort.Strings   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  0runtime.morestack_noctxt   P�  "".autotmp_0564 �Ptype.map.iter[string][]go/token.Position "".path �type.string "".all �type.[]string "".~r2 @Ftype.map[string][]go/token.Position "".~r1 type.[]string "".m  Ftype.map[string][]go/token.Position  ����g�
 � 4�9QhN"?M
  gV�M)? Tgclocals·9f4747e6338c5bdd4db417363b8a0d83 Tgclocals·8744fb04fbd6f74dba2601338d86fe97   :$GOROOT/src/go/build/build.go�"".Import  �  �dH�%    H;a��   H��H1�H��$�   H��$�   H�    H�$H�\$PH�\$H�\$XH�\$H�\$`H�\$H�\$hH�\$ H�\$pH�\$(�    H�T$0H�L$8H�D$@H�T$xH��$�   H��$�   H��H��    �b�����
      X  "".Default   �  ("".(*Context).Import   �  0runtime.morestack_noctxt   ��  
"".~r4 `type.error "".~r3 P type.*"".Package "".mode @$type."".ImportMode "".srcDir  type.string "".path  type.string �|� � �)k 
 f: Tgclocals·5998daf4e6d23f69cd931cd9519af48e Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�"".ImportDir  �  �dH�%    H;avaH��81�H�\$`H�\$hH�    H�$H�\$@H�\$H�\$HH�\$H�\$PH�\$�    H�T$ H�L$(H�D$0H�T$XH�L$`H�D$hH��8��    ����������
      D  "".Default   �  ."".(*Context).ImportDir   �  0runtime.morestack_noctxt   `p  "".~r3 @type.error "".~r2 0 type.*"".Package "".mode  $type."".ImportMode "".dir  type.string p\o � �Q 
 H8 Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�2"".(*Context).shouldBuild  �  �dH�%    H��$X���H;A�8  H��(  H�D$@    H��$8  H��$�   H��$@  H��$H  H��$�   H�� �]  H��$�   H��$�   H��$�   H��$�   H�$H��$�   H�t$H��$�   H�D$�D$
�    L��$�   H��$�   L��$�   H��$�   H��$�   H�D$ H�� �5  H9��%  I��H��L��H��H��H��I��H9��   H)�I)�M��I�� tM�I��L��$�   H��L��$�   H��$�   L��$�   L��$�   L�$H��$�   H�\$H��$�   H�t$�    H��$�   H�l$H��$�   H�L$ H�T$(H��$�   H��$�   H�� �  H��$@  H)�H�\$@H�� �����H�\$@H��$H  H9���  H��H��$8  H��$�   H��$@  H��$�   H��$H  H��$�   �D$?H��$�   H�� ��  H��$�   H��$�   H��$�   H��$�   H�$H��$�   H�L$H��$�   H�D$�D$
�    L��$�   H��$�   L��$�   H��$�   H��$�   H�D$ H�� ��  H9���  I��H��L��H��H��H��I��H9���  H)�I)�M��I�� tM�I��L��$�   H��L��$�   H��$�   L��$�   L��$�   L�$H��$�   H�\$H��$�   H�t$�    H�T$H�L$ H�D$(H��$�   H�$H��$�   H�L$H��$�   H�D$H�    H�\$H�    H�\$ H�    H�\$(�    �\$0�� ��  H�    H��$�   L��$�   H9���  L��$�   H)�I)�I�� tM�L��$  L�$H��$  H�l$L��$   L�D$�    H�L$H�D$ H�l$(H�� �5  H�� �0  ���+�  H�$    H��$�   H�L$H��$�   H�D$H��$�   H�l$�    H�\$ H�H�$H�KH�L$�    H�L$H�D$H�\$ H��$�   H��H��$�   H�� H��$�   ��  H�	H�L$pH�CH�D$xH���I���H�$H�D$H�-    H�l$H�D$   �    �\$ �� �����D$> H��$�   H��$�   H���$  H��H��L��$�   H�� tI��L��$�   H��$   H��$  H��$�   1�H��$�   H�\$HL��$�   L��H�l$HH9���   H�D$XH�� ��   H�H�hH�L$PH�T$pH�l$xH��$0  H�$H�T$`H�T$H�l$hH�l$H��$P  H�\$�    �\$ �� tZ�D$>H�D$XH�L$PH��H��H�l$HH9��{����|$> �	����D$? H��$�   H�� �����\$?��$X  H��(  �멉 �K����    �    ������    �    �����    �    H��I��H9�w0H)�I)�M��I�� tM�	H��$�   L��$�   L��$�   �W����    �    H�,$H�L$H�T$H�    H�\$H�    H�\$ H�    H�\$(�    H��$�   �\$0�� u�����P����    �    H��I��H9�w0H)�I)�M��I�� tM�	H��$�   L��$�   L��$�   ������    �    �������@
      �  bytes.IndexByte   �  bytes.TrimSpace   �	  bytes.IndexByte   �  bytes.TrimSpace   �  "".slashslash   � "".slashslash   �  "".slashslash   �  bytes.HasPrefix   � "".slashslash   �  bytes.TrimSpace   �  2runtime.slicebytetostring   �  strings.Fields   �  $go.string."+build"   �   runtime.eqstring   �  &"".(*Context).match   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  "".slashslash   � "".slashslash   �  "".slashslash   �  bytes.HasPrefix   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   `�  B"".autotmp_0597  type.string "".autotmp_0596 �type.*string "".autotmp_0595  type.int "".autotmp_0594  type.int "".autotmp_0593 �type.string "".autotmp_0591 �type.[]string "".autotmp_0590 _type.[]string "".autotmp_0589  type.int "".autotmp_0588  type.[]uint8 "".autotmp_0587  type.int "".autotmp_0586  type.bool "".autotmp_0585  type.int "".autotmp_0584  type.[]uint8 "".autotmp_0583  type.int "".autotmp_0582  type.[]uint8 "".autotmp_0581  type.int "".autotmp_0578 �type.int "".autotmp_0577  type.int "".autotmp_0576  type.int "".autotmp_0575 /type.[]uint8 "".autotmp_0574 �type.int "".tok �type.string 
"".ok �type.bool "".f �type.[]string "".line �type.[]uint8 "".allok �type.bool "".line �type.[]uint8 "".p �type.[]uint8 "".end �type.int "".~r2 Ptype.bool "".allTags @(type.map[string]bool "".content type.[]uint8 "".ctxt   type.*"".Context ""������ � ��"	(
g`R
 0g`:]r ei�<
)86I
6 @ ����^q��r	�!] Tgclocals·689482aa6db86c01fa54c72fbbe58e52 Tgclocals·6c1e86c4f55eb0f4f23b9aeed94efe32   :$GOROOT/src/go/build/build.go�*"".(*Context).saveCgo  �j  �jdH�%    H��$8���H;A�x  H��H  1�H��$x  H��$�  H��$p  H�$�    H�L$H�D$H��$�   H�$H��$�   H�D$H�    H�\$H�D$   �    H�T$ H�D$(H�L$0H��$�  H��$   H��$  H��$�  1�H��$�  H�D$PH��$�  H��H�l$PH9��8  H��$�   H�� ��  H�H�hH�L$XH��$  H��$  H��$�   H��$�   H��$�   H�$H��$�   H�l$�    H�T$H�L$H����   H��$�   H���*  H��$�   H��   H��uH��$  H�$H��$  H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� t2H��H����  H����� tUH��H����  H�����	t<H��$�   H�L$XH��H��H�l$PH9������1�H��$x  H��$�  H��H  �H��H���8  H��H��H�� tH��H��$8  H�,$H��$@  H�\$�    H�L$H�D$H��$�   H�$H��$�   H�D$H�    H�\$H�D$   �    H��$�   H��$�   H�D$ H�� ��  H��$X  H��$(  H��$`  H��$0  H��$�   H��$  H��$�   H��$   1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �e  HǄ$�     HǄ$�     H��$�  H�    H�$H��$(  H�\$H�D$    �    H�L$H�D$ H��$�  H��$�   H�H��$   �=     ��   H�CH�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$�   H�H��$   �=     ufH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$x  H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H9���  H��H��H��H��H��H9���  H)�I��H�� tM�L��$H  H��$P  H��$�   H�$H��$�   H�t$�    L�L$L��$h  H�D$H�T$ H��$x  H��$p  H����  H��$X  H��$(  H��$`  H��$0  H��$�   H��$  H��$�   H��$   1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �e  HǄ$�     HǄ$�     H��$�  H�    H�$H��$(  H�\$H�D$    �    H�L$H�D$ H��$�  H��$�   H�H��$   �=     ��   H�CH�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$�   H�H��$   �=     ufH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$x  H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H��H��H9��9  H��H��H��L��H9��  H��H�H�L�CL��$�  H��$�  H��$8  H��$�   L��$@  L��$�   H��$�  H�� ��   1�@�t$GH��$�  1�H��$�  H�|$`L��$�  L��H�l$`H9�}|H��H�D$xH�� ��  H� H�kH�L$hH��$8  H��$@  H��$P  H�$H��$�   H�D$H��$�   H�l$H�D$    �    �t$G�\$ �� �  H��   @�� �����H��$H  H�$H��$P  H�\$�    H�l$H��$  H�T$H��$  H�L$ H��$   H�D$(H�\$0H��$�   H��$�   H�� ��  H��$X  H��$(  H��$`  H��$0  H��$�   H��$  H��$�   H��$   1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �e  HǄ$�     HǄ$�     H��$�  H�    H�$H��$(  H�\$H�D$    �    H�L$H�D$ H��$�  H��$�   H�H��$   �=     ��   H�CH�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$�   H�H��$   �=     ufH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$x  H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H��$�  1�H��$�  H�T$hH��$�  H��H�l$hH9���  H��H�L$xH�� �e  H�	H�kH�D$pH�D$HH��$8  H��$@  H��$X  H�$H��$`  H�l$H��$h  H�|$H�H�H�NH�O�    H�T$ H�L$(�\$0�� ��  H��$X  H��$  H��$`  H��$   H��$X  H��$(  H��$`  H��$0  1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �e  HǄ$�     HǄ$�     H��$�  H�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��$�   H�H��$   �=     ��   H�CH�    H�$H��$(  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$�   H�H��$   �=     ufH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$x  H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H��$  H�l$HL��$  L9���  H��H�H��$`  H�KH��$X  �=     ��  H�H�L$xH�D$pH��H��H�l$hH9��4���H��$�   H��$8  H��$�   H��|TH���@  H�$H��$@  H�D$H�-    H�l$H�D$   �    H��$8  H��$@  H�\$ H�� ��  H���	  H�$H��$@  H�D$H�-    H�l$H�D$   �    L��$  H��$8  H��$@  �\$ �� ��  H��$h  H�� ��  H��   H��  H��  H��$�  H��$�  H��$�  H��H��$�  L�H)�H�� ~[H�    H�$H��$�  H�t$H�|$H��$�  H�D$H�L$ �    L��$  H��$�  H�t$(H�\$0H��$�  H�D$8H�    H�$H��H��L�I��H��$�  H9���   H9���   H)�I)�I��H��$�  I�� tHk�I�H�l$L�D$L�L$H��$  H�\$ L�T$(H��$   H�\$0�    H��$�  H��$�  H��$  H�H9�wPH��H��$h  H��  H��  H��$�  �=     uH��   ����L��   L�$H�l$�    ������    �    ��Z���H��$@  H����  H�$H�D$H�-    H�l$H�D$   �    L��$  �\$ �� ��  H��$h  H�� ��  H��H  H��P  H��X  H��$�  H��$�  H��$�  H��H��$�  L�H)�H�� ~[H�    H�$H��$�  H�t$H�T$H��$�  H�D$H�L$ �    L��$  H��$�  H�t$(H�\$0H��$�  H�D$8H�    H�$H��H��L�I��H��$�  H9���   H9���   H)�I)�I��H��$�  I�� tHk�I�H�l$L�D$L�L$H��$  H�\$ L�T$(H��$   H�\$0�    H��$�  H��$�  H��$  H�H9�wPH��H��$h  H��P  H��X  H��$�  �=     uH��H  ����L��H  L�$H�l$�    ������    �    ��Z���H��$X  H��$  H��$`  H��$   H��$�   H��$(  H��$�   H��$0  1�H��$(  H��$0  H��$8  H��$@  H��$(  H�� �e  HǄ$�     HǄ$�     H��$�  H�    H�$H��$  H�\$H�D$    �    H�L$H�D$ H��$�  H��$�   H�H��$   �=     ��   H�CH�    H�$H��$(  H�\$H�D$    �    H�L$H�D$ H��$�  H��H��$�   H�H��$   �=     ufH�CH�    H�$H�D$   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�L$(H�D$0H��$x  H��$�  H��H  �L�CL�$H�D$�    �L�CL�$H�D$�    ���������H���	  H�$H��$@  H�D$H�-    H�l$H�D$   �    L��$  H��$8  H��$@  �\$ �� ��  H��$h  H�� ��  H��  H��   H��(  H��$�  H��$�  H��$�  H��H��$�  L�H)�H�� ~[H�    H�$H��$�  H�t$H�T$H��$�  H�D$H�L$ �    L��$  H��$�  H�t$(H�\$0H��$�  H�D$8H�    H�$H��H��L�I��H��$�  H9���   H9���   H)�I)�I��H��$�  I�� tHk�I�H�l$L�D$L�L$H��$  H�\$ L�T$(H��$   H�\$0�    H��$�  H��$�  H��$  H�H9�wPH��H��$h  H��   H��(  H��$�  �=     uH��  ����L��  L�$H�l$�    �����    �    ��Z���H���	  H�$H��$@  H�D$H�-    H�l$H�D$   �    L��$  H��$8  H��$@  �\$ �� ��  H��$h  H�� ��  H��0  H��8  H��@  H��$�  H��$�  H��$�  H��H��$�  L�H)�H�� ~[H�    H�$H��$�  H�t$H�|$H��$�  H�D$H�L$ �    L��$  H��$�  H�t$(H�\$0H��$�  H�D$8H�    H�$H��H��L�I��H��$�  H9���   H9���   H)�I)�I��H��$�  I�� tHk�I�H�l$L�D$L�L$H��$  H�\$ L�T$(H��$   H�\$0�    H��$�  H��$�  H��$  H�H9�wPH��H��$h  H��8  H��@  H��$�  �=     uH��0  ����L��0  L�$H�l$�    ������    �    ��Z���H��$@  H��
�����H�$H�D$H�-    H�l$H�D$
   �    L��$  �\$ �� �����H��$h  H�� ��  H��`  H��h  H��p  H��$�  H��$�  H��$�  H��H��$�  L�H)�H�� ~[H�    H�$H��$�  H�t$H�|$H��$�  H�D$H�L$ �    L��$  H��$�  H�t$(H�\$0H��$�  H�D$8H�    H�$H��H��L�I��H��$�  H9���   H9���   H)�I)�I��H��$�  I�� tHk�I�H�l$L�D$L�L$H��$  H�\$ L�T$(H��$   H�\$0�    H��$�  H��$�  H��$  H�H9�wPH��H��$h  H��h  H��p  H��$�  �=     uH��`  ����L��`  L�$H�l$�    ������    �    ��Z���H�$H�T$�    �=����    �����H�D$xH�L$hH��H���c���� �x����    �    �    �    �    �    �    �    � �X����    �c�����̀
      �  6go/ast.(*CommentGroup).Text   �  go.string."\n"   �  strings.Split   �  "strings.TrimSpace   �   go.string."#cgo"   �   runtime.eqstring   �	  "strings.TrimSpace   �
  go.string.":"   �
  strings.Index   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  Jgo.string."%s: invalid #cgo line: %s"   �  fmt.Errorf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  strings.Fields   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  Jgo.string."%s: invalid #cgo line: %s"   �  fmt.Errorf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �   &"".(*Context).match   �!  "".splitQuoted   �%  type.string   �%  runtime.convT2E   �& (runtime.writeBarrier   �&  type.string   �&  runtime.convT2E   �' (runtime.writeBarrier   �'  Jgo.string."%s: invalid #cgo line: %s"   �(  fmt.Errorf   �)  .runtime.writebarrierptr   �)  .runtime.writebarrierptr   �,  "".expandSrcDir   �/  type.string   �/  runtime.convT2E   �0 (runtime.writeBarrier   �0  type.string   �1  runtime.convT2E   �1 (runtime.writeBarrier   �2  Vgo.string."%s: malformed #cgo argument: %s"   �3  fmt.Errorf   �3  .runtime.writebarrierptr   �4  .runtime.writebarrierptr   �5 (runtime.writeBarrier   �7  &go.string."LDFLAGS"   �7  "runtime.cmpstring   �8  $go.string."CFLAGS"   �8   runtime.eqstring   �:  type.[]string   �;  &runtime.growslice_n   �<  type.string   �>  ,runtime.typedslicecopy   �? (runtime.writeBarrier   �?  .runtime.writebarrierptr   �?  $runtime.panicslice   �?  $runtime.panicslice   �@  &go.string."LDFLAGS"   �@   runtime.eqstring   �B  type.[]string   �C  &runtime.growslice_n   �D  type.string   �F  ,runtime.typedslicecopy   �G (runtime.writeBarrier   �G  .runtime.writebarrierptr   �G  $runtime.panicslice   �H  $runtime.panicslice   �J  type.string   �K  runtime.convT2E   �K (runtime.writeBarrier   �L  type.string   �L  runtime.convT2E   �M (runtime.writeBarrier   �M  Jgo.string."%s: invalid #cgo verb: %s"   �N  fmt.Errorf   �O  .runtime.writebarrierptr   �O  .runtime.writebarrierptr   �P  (go.string."CPPFLAGS"   �P   runtime.eqstring   �R  type.[]string   �S  &runtime.growslice_n   �S  type.string   �U  ,runtime.typedslicecopy   �V (runtime.writeBarrier   �W  .runtime.writebarrierptr   �W  $runtime.panicslice   �W  $runtime.panicslice   �X  (go.string."CXXFLAGS"   �X   runtime.eqstring   �Z  type.[]string   �[  &runtime.growslice_n   �\  type.string   �^  ,runtime.typedslicecopy   �_ (runtime.writeBarrier   �_  .runtime.writebarrierptr   �_  $runtime.panicslice   �`  $runtime.panicslice   �`  ,go.string."pkg-config"   �a   runtime.eqstring   �b  type.[]string   �c  &runtime.growslice_n   �d  type.string   �f  ,runtime.typedslicecopy   �g (runtime.writeBarrier   �g  .runtime.writebarrierptr   �h  $runtime.panicslice   �h  $runtime.panicslice   �h  .runtime.writebarrierptr   �h  $runtime.panicindex   �i  $runtime.panicindex   �i  $runtime.panicslice   �i  $runtime.panicslice   �i  $runtime.panicslice   �i  $runtime.panicslice   �i  $runtime.panicindex   �i  $runtime.panicindex   �j  $runtime.panicslice   �j  0runtime.morestack_noctxt   p�	  �"".autotmp_0689  "type.interface {} "".autotmp_0688  "type.interface {} "".autotmp_0687  (type.[2]interface {} "".autotmp_0685  *type.*[2]interface {} "".autotmp_0684  &type.[]interface {} "".autotmp_0683  type.int "".autotmp_0682  type.[]string "".autotmp_0681  type.[]string "".autotmp_0680  type.int "".autotmp_0679  type.[]string "".autotmp_0678  type.[]string "".autotmp_0677  type.int "".autotmp_0676  type.[]string "".autotmp_0675  type.[]string "".autotmp_0674  type.int "".autotmp_0673  type.[]string "".autotmp_0672  type.[]string "".autotmp_0671  type.int "".autotmp_0670 �type.[]string "".autotmp_0669  type.[]string "".autotmp_0668  type.string "".autotmp_0667  "type.interface {} "".autotmp_0666  "type.interface {} "".autotmp_0665  (type.[2]interface {} "".autotmp_0663  *type.*[2]interface {} "".autotmp_0662  &type.[]interface {} "".autotmp_0661  type.string "".autotmp_0660  type.*string "".autotmp_0659  type.int "".autotmp_0658  type.int "".autotmp_0657  "type.interface {} "".autotmp_0656  "type.interface {} "".autotmp_0655  (type.[2]interface {} "".autotmp_0653  *type.*[2]interface {} "".autotmp_0652  &type.[]interface {} "".autotmp_0651  type.string "".autotmp_0650 �type.*string "".autotmp_0649  type.int "".autotmp_0648  type.int "".autotmp_0647  type.string "".autotmp_0645  "type.interface {} "".autotmp_0644  "type.interface {} "".autotmp_0643  (type.[2]interface {} "".autotmp_0641  *type.*[2]interface {} "".autotmp_0640  &type.[]interface {} "".autotmp_0639  "type.interface {} "".autotmp_0638 �"type.interface {} "".autotmp_0637 ?(type.[2]interface {} "".autotmp_0634 �&type.[]interface {} "".autotmp_0633 �type.string "".autotmp_0632 �type.*string "".autotmp_0631 �type.int "".autotmp_0630 �type.int "".autotmp_0629  type.error "".autotmp_0628  type.string "".autotmp_0627  type.string "".autotmp_0626  type.error "".autotmp_0625  type.string "".autotmp_0624  type.string "".autotmp_0623  type.[]string "".autotmp_0622  type.error "".autotmp_0621  type.string "".autotmp_0620  type.string "".autotmp_0618  type.[]string "".autotmp_0617  type.int "".autotmp_0616 �type.int "".autotmp_0615 �type.[]string "".autotmp_0614 �type.int "".autotmp_0613  type.int "".autotmp_0612  type.error "".autotmp_0611  type.string "".autotmp_0610  type.string "".autotmp_0609  type.int "".autotmp_0607  type.int "".autotmp_0606  type.string "".autotmp_0604 �type.string "".autotmp_0603 �type.string "".autotmp_0602 �type.string "".autotmp_0601  type.string "".autotmp_0600 �type.int "".autotmp_0599 �type.[]string "".autotmp_0598 �type.[]string "".arg �type.string "".i �type.int "".err �type.error "".args otype.[]string "".c �type.string 
"".ok �type.bool "".verb �type.string "".cond �type.[]string "".f �type.[]string "".argstr �type.string "".line �type.string "".orig �type.string "".line �type.string "".text �type.string "".~r3 Ptype.error 
"".cg @2type.*go/ast.CommentGroup 
"".di 0 type.*"".Package "".filename type.string "".ctxt   type.*"".Context h"�	��	�	��	�	��	�	��	�	��	�	��	�	��	 �5 ��4�
(�"�kFH
�A=�bZG

W�cQ�Ir[�ijij
K�uvuv�[�mnmn[�qrqrK�yzyz		 � @�n�=��4��4�B��4�
�	�4���k
E��k
��4U��k
E��k
E��k

w Tgclocals·5f7cd344685fbb4cd325c2c2d65d66f9 Tgclocals·456125ec998d6bb6d5850305cab89579   :$GOROOT/src/go/build/build.go�"".expandSrcDir  �  �dH�%    H�D$�H;A��  H��   1�H��$�   H��$�   H��$�   H�$H��$�   H�\$�    H�\$H��$�   H�\$H��$�   H��$�   H�$H��$�   H�\$H�    H�\$H�D$	   �    H�\$ H�\$xH�\$(H��$�   H�\$0H��$�   H��$�   H��}ZH��$�   H�$H��$�   H�\$�D$ �    �\$H��H��$�   H��$�   H��$�   H��$�   ��$�   H�Ĩ   �H��   H�T$xH��$�   H��$�   H��$�   1�H��$�   H�L$@H��$�   H�l$@H9�}wH�T$PH�� �V  H�:H�JH�t$HH�|$hH�|$XH�L$pH�L$`< �'  H�� �  H�<$H�L$�D$ �    H�t$HH�T$P�\$H��H��H��H�l$@H9�|�< ��   H��$�   H�� ��   H��$�   H�$H��$�   H�\$�D$�    �\$�\$?H�\$xH�$H��$�   H�\$H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�L$(H�D$0H��$�   H��$�   �|$? tH�� ��$�   H�Ĩ   �Ƅ$�    ���D$?�u����D$? �k���H��   ����1�����������    �����������������
      �  *path/filepath.ToSlash   �  *go.string."${SRCDIR}"   �  strings.Split   �  "".safeCgoName   �  "".safeCgoName   �  "".safeCgoName   �	  strings.Join   �  0runtime.morestack_noctxt   p�  "".autotmp_0698 type.string "".autotmp_0697 �type.*string "".autotmp_0696 �type.int "".autotmp_0695  type.int "".autotmp_0694  type.bool "".autotmp_0693  type.bool "".autotmp_0692 /type.[]string "".autotmp_0690 �type.int "".chunk �type.string 
"".ok �type.bool "".chunks _type.[]string "".~r3 `type.bool "".~r2 @type.string "".srcdir  type.string "".str  type.string .�������8� � D�18WZm7FL5  J�`K� Tgclocals·776d9d553b2634d9ea530b3c76543df4 Tgclocals·6347b58243cc1c5f8f735d259ec00f70   :$GOROOT/src/go/build/build.go�"".safeCgoName  �  �dH�%    H;a�  H��HH�T$XH�� u
�D$h H��H�H�    H�\$0H�    H�\$8H�    H�\$@�|$` u7H�\$8H�l$@H����   H��H��L�D$0H�� tI��H�\$8H�l$@L�D$01�H9�}jH�\$PH�L$(H9�seH��+@���sFH�\$0H�$H�\$8H�\$H�\$@H�\$@�l$�    H�T$XH�L$(H�\$ H�� }
�D$h H��H�H��H9�|��D$hH��H��    �    �    ��������������������
      ^  "".safeBytes   v "".safeBytes   �  "".safeBytes   �  bytes.IndexByte   �  $runtime.panicindex   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0699  type.int "".i ?type.int "".safe /type.[]uint8 "".~r2 0type.bool "".spaces  type.bool "".s  type.string 8��������� � <�
$7X


  �6' Tgclocals·f47057354ec566066f8688a4970cff5a Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60   :$GOROOT/src/go/build/build.go�"".splitQuoted  �  �dH�%    H��$h���H;A�q  H��  1�1�1�H��$H  H��$P  1�H��$0  H��$8  H��$@  1�H��$�   H��$�   H��$�   H��$(  H�    H�$H�D$H�D$�    H�\$H��$   H�\$ H��$  H�\$(H��$  �D$G �D$F �D$L    H�D$P    H��$   H��$�   H��$(  H��$�   H�D$`    H�\$`H�\$XH��$�   H�$H��$�   H�\$H�\$`H�\$�    H��$   �t$LH�L$PH�\$H�\$`�D$ H�\$`H�� ��  �|$G t/�D$G L��$  L9�sH���H��H��H�\$P�q����    ��\u
�D$G�[����� t9�u��D$L    �E�����"�|  ��'�s  �D$H�$�    H��$   H�L$P�D$H�\$�� �t����|$F u
H�� ������D$F H��$  H9��  H�$    H��$�   H�|$H��$�   H�L$H��$�   H�l$�    H�\$ H��$�   H�\$(H��$�   H��$�   H��$�   H��$�   H��H��H9�wSH��$�   H��H��Hk�H�H��$�   H�kH��$�   �=     uH�+H�D$P    �-���H�$H�l$�    ��H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�   H��$�   H��$�   �_����    �D$F�D$L�����|$F �  H�� ��  �� �  H�    H��$�   HǄ$�      1�H��$�   H��$�   H�    H�$�    H�D$H�D$hH��$�   H�hH��$�   �=     ��   H�(H�D$hH�    1�H9�tMH�L$hH��$H  H��$P  H��$�   H��$0  H��$�   H��$8  H��$�   H��$@  H��  �H�    H�$H�    H�\$H�    H�\$�    H�D$�H�$H�l$�    H�D$h�Y����|$G �v���H�    H��$�   HǄ$�      1�H�\$pH�\$xH�    H�$�    H�D$H�D$hH��$�   H�hH��$�   �=     u_H�(H�D$hH�    1�H9�tH�T$hH��$H  H��$P  �����H�    H�$H�    H�\$H�    H�\$�    H�D$�H�$H�l$�    H�D$h�H��$  H9��   H�$    H��$�   H�|$H��$�   H�L$H��$�   H�l$�    �t$LH�\$ H��$�   H�\$(H��$�   H��$�   H��$�   H��$�   H��H��H9�wQH��$�   H��H��Hk�H�H��$�   H�kH��$�   �=     uH�+�H���H�$H�l$�    �t$L�1���H�-    H�,$H�L$H�D$H�T$H�\$ �    �t$LH�L$(H�\$0H�T$8H��H��H��$�   H��$�   H��$�   �]����    �    �j�������������N
      �  type.[]int32   �  "runtime.makeslice   �  &runtime.stringiter2   �  $runtime.panicindex   �  unicode.IsSpace   �	  2runtime.slicerunetostring   �
 (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  $runtime.panicslice   �  4go.string."unclosed quote"   �  .type.errors.errorString   �  "runtime.newobject   � (runtime.writeBarrier   �  Bgo.itab.*errors.errorString.error   �  0type.*errors.errorString   �  type.error   �  Bgo.itab.*errors.errorString.error   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  >go.string."unfinished escaping"   �  .type.errors.errorString   �  "runtime.newobject   � (runtime.writeBarrier   �  Bgo.itab.*errors.errorString.error   �  0type.*errors.errorString   �  type.error   �  Bgo.itab.*errors.errorString.error   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  2runtime.slicerunetostring   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   p�  :"".autotmp_0720  type.*uint8 "".autotmp_0719  type.error "".autotmp_0718  0type.*errors.errorString "".autotmp_0715 �0type.*errors.errorString "".autotmp_0714  type.string "".autotmp_0713 �type.string "".autotmp_0711  type.int "".autotmp_0710 �type.int "".autotmp_0709  0type.*errors.errorString "".autotmp_0708  0type.*errors.errorString "".autotmp_0707  type.[]int32 "".autotmp_0706  type.int "".autotmp_0705 �type.[]int32 "".autotmp_0703 �type.string "".autotmp_0702 �type.int "".~r0 �type.error errors.text·2 �type.string "".~r0 �type.error errors.text·2 �type.string "".rune �type.int32 "".i �type.int "".quote �type.int32 "".quoted �type.bool "".escaped �type.bool "".arg /type.[]int32 "".args _type.[]string "".err Ptype.error "".r  type.[]string "".s  type.string ""������ � ��RI	�*10'	+�	'&]6	�8G�D	�aE D ��bE�7k
�aa	�; Tgclocals·80238e4f21dcc74d0e33ebfc08caa30e Tgclocals·3766546ec9671d5836402e8fa0c9f6e2   :$GOROOT/src/go/build/build.go�&"".(*Context).match  �$  �$dH�%    H�D$�H;A��  H���   H��$  H��$�   H��$   H�� uX1�H9�tAH��$�   H��$�   �D$+H�    H�$H�T$H��$�   H�\$H�\$+H�\$�    Ƅ$   H���   �H�$H�D$H�    H�\$H�D$   �    L��$  H��$�   H��$   H�D$ H�� ��   H�D$0H9���   H��$�   H�$H��$�   H�|$H��$�   H�D$L�T$�    �\$ �\$*H�\$0H��H��$   H9�wrL��$�   H)�H�� tM�H��$�   H�$L��$�   L�D$H��$�   H�l$H��$  H�\$�    �\$ �|$* t��$  H���   �Ƅ$   ���    �    H��$�   L�    L��$�   H��   H��$�   H��$�   H9��  H9��  H9���  H��$�   H�<$H��$�   H�D$L�D$H�D$�    L��$  H��$�   H��$   �\$ H��< tƄ$   H���   �H�|$pL�    L��$�   H��   H�L$xH��$�   H9��]  H9��M  H9��=  H��$�   H�<$H��$�   H�D$L�D$H�D$�    L��$  H��$�   H��$   �\$ H��< t}H��~mH��H��r]H��H��H�� tH��H��H��$�   H�$H��$�   H�l$H��$�   H�L$L�T$�    �\$ H��H����$  H���   ��    Ƅ$   ��1�I9�tQH��$�   H��$�   �D$+H�    H�$L�T$H��$�   H�\$H�\$+H�\$�    H��$�   H��$   H��$�   H��$�   1�H�T$@H��$�   H�$H��$�   H�\$H�T$�    H��$   H�T$�D$ H�T$8H�� tY�D$,�$�    H�T$8�\$�� u9�\$,�$�    H�T$8�L$,�\$�� u��_t��.tƄ$   H���   ��c���H��$�   �]@�� tSH��uMH��$�   H�,$H�L$H�-    H�l$H�D$   �    H��$   �\$ �� tƄ$  H���   �H��$�   H�� ��  H�SH�CH9�uRH��$�   H�,$H�L$H��$�   H�T$H��$�   H�D$�    H��$   �\$ �� tƄ$  H���   �H��$�   H�� �x  H�H�CH9�uBH��$�   H�,$H�L$H��$�   H�T$H��$�   H�D$�    H��$   �\$ �� u�H��$�   H�� �  H�SHH�CPH9�uFH��$�   H�,$H�L$H��$�   H�T$H��$�   H�D$�    H��$   �\$ �� �+���H��$�   H�� ��  H�SH�CH����   H��$�   H�$H��$�   H�D$H�-    H�l$H�D$   �    H��$   �\$ �� tSH��uMH��$�   H�,$H�L$H�-    H�l$H�D$   �    H��$   �\$ �� tƄ$  H���   �H��$�   H�� ��  H�SXH�C`H�khH��$�   1�H��$�   H�D$@H��$�   H�l$@H9���   H�T$HH�� ��  H�:H�BH�t$8H��$�   H�|$`H��$�   H�D$hH9�uLH�<$H�D$H��$�   H�l$H�L$�    H�t$8H�T$HH��$   �\$ �� tƄ$  H���   �H��H��H�l$@H9��e���H��$�   H�� ��   H�SpH�CxH���   H��$�   1�H��$�   H�D$@H��$�   H�l$@H9���   H�T$HH�� ��   H�:H�BH�t$8H��$�   H��$�   H9�uVH�|$PH�<$H�D$XH�D$H��$�   H�l$H�L$�    H�t$8H�T$HH��$   �\$ �� tƄ$  H���   �H��H��H�l$@H9��e���Ƅ$   H���   É�]����������f����������T����������������	���1������    1������1��P����    1��B����    �����������������D
      �  (type.map[string]bool   �  $runtime.mapassign1   �  go.string.","   �  strings.Index   �  &"".(*Context).match   �  &"".(*Context).match   �  $runtime.panicslice   �  $runtime.panicslice   �  go.string."!!"   �   runtime.eqstring   �	  go.string."!"   �   runtime.eqstring   �  &"".(*Context).match   �  $runtime.panicslice   �  (type.map[string]bool   �  $runtime.mapassign1   �  &runtime.stringiter2   �   unicode.IsLetter   �  unicode.IsDigit   �  go.string."cgo"   �   runtime.eqstring   �   runtime.eqstring   �   runtime.eqstring   �   runtime.eqstring   �  &go.string."android"   �   runtime.eqstring   �  "go.string."linux"   �   runtime.eqstring   �   runtime.eqstring   �!   runtime.eqstring   �#  $runtime.panicslice   �#  $runtime.panicslice   �$  0runtime.morestack_noctxt   P�  b"".autotmp_0768  type.string "".autotmp_0767  type.*string "".autotmp_0766  type.int "".autotmp_0765  type.int "".autotmp_0764  type.string "".autotmp_0763 �type.*string "".autotmp_0762  type.int "".autotmp_0761  type.int "".autotmp_0760  type.string "".autotmp_0759  type.string "".autotmp_0758  type.string "".autotmp_0757  type.string "".autotmp_0755  type.int "".autotmp_0754  type.int "".autotmp_0753  type.bool "".autotmp_0751  type.[]string "".autotmp_0750 /type.[]string "".autotmp_0748  type.bool "".autotmp_0747  type.string "".autotmp_0746  type.bool "".autotmp_0745  type.string "".autotmp_0744  type.bool "".autotmp_0743  type.string "".autotmp_0742  type.int "".autotmp_0741  type.string "".autotmp_0740  type.int "".autotmp_0739  type.int "".autotmp_0738  type.int "".autotmp_0737  type.string "".autotmp_0736 �type.int "".autotmp_0734  type.int "".autotmp_0733  type.string "".autotmp_0732 �type.int "".autotmp_0731 otype.string "".autotmp_0730 �type.bool "".autotmp_0729 Otype.string "strings.prefix·3 �type.string strings.s·2 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "".tag �type.string "".tag �type.string "".c �type.int32 "".ok1 �type.bool "".i �type.int "".~r2 @type.bool "".allTags 0(type.map[string]bool "".name type.string "".ctxt   type.*"".Context ��u��������������h��p�����������$��b� � ��7AJGg ��}Q
VDTa��{F
yK		' , �3�J���9 Tgclocals·a4a72fe4111c0d730d77d6113711d8c8 Tgclocals·a95d0301643df1b330639fcf326ec36f   :$GOROOT/src/go/build/build.go�8"".(*Context).goodOSArchFile  �&  �&dH�%    H�D$�H;A�u	  H��   H��$�   H�$H��$�   H�\$H�    H�\$H�D$   �    H��$�   H�D$ H���tH9��	  H��H��$�   H�$H��$�   H�L$H�    H�\$H�D$   �    H�D$ H�� }Ƅ$�   H�Ĉ   �H��$�   H9���  L��$�   H)�H�� tM� L��$�   L�$H��$�   H�l$H�    H�\$H�D$   �    H�\$ H�\$pH�T$(H�\$0H��$�   H�� ��   H��H�T$HH��H�l$pH�T$xH9��  H��H�H�M H�L$`H�EH�D$hH��uNH�$H�D$H�-    H�l$H�D$   �    H�T$x�\$ �� tH�\$HH��H��$�   H9���  H��H��H����  H�    H�$H�    H�\$H��H�D$@H�t$pH��H�T$xH9��^  H��H�H�|$H�H�H�NH�O�    H�T$xH�D$@H�\$ �+@�� �>  H�    H�$H�    H�\$H��H��H�t$pH9���  H��H�H�|$H�H�H�NH�O�    H��$�   H�T$xH�D$@H�\$ �+@�� ��  1�H9���   �D$?H��H��H�    H�$H�t$H�\$pH9���  H��H�H�\$H�\$?H�\$�    �D$?H�l$@H��H�    H�$H��$�   H�\$H�\$pL�D$xL9��:  H��H�H�\$H�\$?H�\$�    H�T$xH�D$@H��H��H�l$pH9���  H��H�H�u H�MH��$�   H�� ��  H�H�CH9���  H�t$`H�4$H�L$hH�L$H�T$PH�T$H�D$XH�D$�    �\$ �� �x  H��$�   H�� �_  H�KH�CH����   H�L$PH�$H�D$XH�D$H�-    H�l$H�D$   �    �\$ �� txH�\$@H�l$pL�D$xH��L9���   H��H�H�M H�EH��uGH�L$PH�$H�D$XH�D$H�-    H�l$H�D$   �    �\$ �� tƄ$�   H�Ĉ   �H�\$@H�l$pL�D$xH��L9�sxH��H�H�U H�EH��$�   H�� tWH�sH�KH9�u@H�T$PH�$H�D$XH�D$H�t$`H�t$H�L$hH�L$�    �\$ ��$�   H�Ĉ   �Ƅ$�    ����    �    �����Ƅ$�    H�Ĉ   É�'����    �    �    H���P  H�    H�$H�    H�\$H��H�D$@H��H�t$pH�T$xH9���  H��H�H�|$H�H�H�NH�O�    H��$�   H�T$xH�D$@H�\$ �+@�� ��  1�H9�tN�D$?H��H��H�    H�$H�t$H�\$pH9���  H��H�H�\$H�\$?H�\$�    H�T$xH�D$@H��$�   H�� �c  H�sH�KH����   H�t$PH�4$H�L$XH�L$H�-    H�l$H�D$   �    H�T$xH�D$@�\$ �� tzH��H��H�l$pH9���   H��H�H�u H�MH��uQH�t$PH�4$H�L$XH�L$H�-    H�l$H�D$   �    H�T$xH�D$@�\$ �� tƄ$�   H�Ĉ   �H��H��H�l$pH9�sxH��H�H�U H�EH��$�   H�� tWH�sH�KH9�u@H�T$PH�$H�D$XH�D$H�t$`H�t$H�L$hH�L$�    �\$ ��$�   H�Ĉ   �Ƅ$�    ����    �    ������    H���\  H�    H�$H�    H�\$H��H�D$@H��H�t$pH�T$xH9��7  H��H�H�|$H�H�H�NH�O�    H��$�   H�\$ �+@�� ��   1�H9�tK�D$?H�l$@H��H�    H�$H�L$H�\$pL�D$xL9���   H��H�H�\$H�\$?H�\$�    H�\$@H��H�l$pL�D$xL9�swH��H�H�u H�MH��$�   H�� tVH�H�CH9�u@H�t$`H�4$H�L$hH�L$H�T$PH�T$H�D$XH�D$�    �\$ ��$�   H�Ĉ   �Ƅ$�    ����    �    Ƅ$�   H�Ĉ   ��    �    �    �    �    �    �    �    �    �i������������x
      v  go.string."."   �  strings.Index   �  go.string."_"   �  strings.Index   �  go.string."_"   �  strings.Split   �   go.string."test"   �   runtime.eqstring   �  (type.map[string]bool   �  "".knownOS   �  4runtime.mapaccess1_faststr   �	  (type.map[string]bool   �	  "".knownArch   �
  4runtime.mapaccess1_faststr   �  (type.map[string]bool   �  $runtime.mapassign1   �  (type.map[string]bool   �  $runtime.mapassign1   �   runtime.eqstring   �  &go.string."android"   �   runtime.eqstring   �  "go.string."linux"   �   runtime.eqstring   �   runtime.eqstring   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  (type.map[string]bool   �  "".knownOS   �  4runtime.mapaccess1_faststr   �  (type.map[string]bool   �  $runtime.mapassign1   �  &go.string."android"   �   runtime.eqstring   �  "go.string."linux"   �   runtime.eqstring   �   runtime.eqstring   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  (type.map[string]bool   �  "".knownArch   �   4runtime.mapaccess1_faststr   �!  (type.map[string]bool   �"  $runtime.mapassign1   �$   runtime.eqstring   �$  $runtime.panicindex   �$  $runtime.panicindex   �%  $runtime.panicindex   �%  $runtime.panicindex   �%  $runtime.panicindex   �%  $runtime.panicindex   �%  $runtime.panicslice   �%  $runtime.panicindex   �&  $runtime.panicslice   �&  $runtime.panicslice   �&  0runtime.morestack_noctxt   P�  <"".autotmp_0794  type.string "".autotmp_0793  type.string "".autotmp_0792  type.int "".autotmp_0791  type.string "".autotmp_0790  type.string "".autotmp_0789  type.string "".autotmp_0788  type.string "".autotmp_0787  type.int "".autotmp_0786  type.string "".autotmp_0785  type.string "".autotmp_0784  type.string "".autotmp_0783  type.string "".autotmp_0782 otype.string "".autotmp_0781  type.string "".autotmp_0780  type.int "".autotmp_0779  type.int "".autotmp_0778 Otype.string "".autotmp_0777  type.bool "".autotmp_0776  type.bool "".autotmp_0775  type.bool "".autotmp_0774  type.bool "".autotmp_0773  type.bool "".autotmp_0772 �type.bool "".n �type.int "".n type.int "".l /type.[]string "".~r2 @type.bool "".allTags 0(type.map[string]bool "".name type.string "".ctxt   type.*"".Context |����������2�����y�����+��8� � ��F8&Oy�E]���N��xK� 0 M������� Tgclocals·c9451ec7b4e00af2b1e38fde82914877 Tgclocals·ac1513c540ef28dcd9fb2a42fdde591a   :$GOROOT/src/go/build/build.go�"".init.1  �	  �	dH�%    H�D$�H;A�  H��   H�    H�$H�D$Q   �    H�T$H�D$H�L$ H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$0H��$�   H��H�l$0H9���   H�D$@H�� ��  H�H�hH�L$8H�T$hH�l$pH�T$HH�T$xH�l$PH��$�   �D$/H�    H�$H�    H�\$H�\$xH�\$H�\$/H�\$�    H�D$@H�L$8H��H��H�l$0H9��p���H�    H�$H�D$�   �    H�T$H�D$H�L$ H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$0H��$�   H��H�l$0H9���   H�D$@H�� ��   H�H�hH�L$8H�T$hH�l$pH�T$XH�T$xH�l$`H��$�   �D$/H�    H�$H�    H�\$H�\$xH�\$H�\$/H�\$�    H�D$@H�L$8H��H��H�l$0H9��p���H�ĸ   É �p���� �i����    ������
      D  �go.string."android darwin dragonfly freebsd linux nacl netbsd openbsd plan9 solaris windows "   h  strings.Fields   �  (type.map[string]bool   �  "".knownOS   �  $runtime.mapassign1   �  ""..gostring.1   �  strings.Fields   �  (type.map[string]bool   �  "".knownArch   �  $runtime.mapassign1   �  0runtime.morestack_noctxt    �  $"".autotmp_0810  type.string "".autotmp_0809  type.*string "".autotmp_0808  type.int "".autotmp_0807  type.int "".autotmp_0806 �type.string "".autotmp_0805 �type.*string "".autotmp_0804 �type.int "".autotmp_0803 �type.int "".autotmp_0802  type.bool "".autotmp_0801  type.string "".autotmp_0800  type.[]string "".autotmp_0799  type.[]string "".autotmp_0798 �type.bool "".autotmp_0797 type.string "".autotmp_0796 _type.[]string "".autotmp_0795 /type.[]string "".v �type.string "".v �type.string  ����� � 4��L�L  3�8�E Tgclocals·69c1753bd5f81501d95132d08af04464 Tgclocals·30fa7c694f0b53328be0204760229368   :$GOROOT/src/go/build/build.go� "".IsLocalImport  �  �dH�%    H;a��  H��xH��$�   H����  H��$�   H�$H�|$H�    H�\$H�D$   �    H��$�   �\$ H��< �x  H���g  H��$�   H�$H�|$H�    H�\$H�D$   �    H��$�   �\$ H��< �  L��$�   L�L$(L�    L�D$HH��   H�|$0H�D$PH9���   H9���   H9���   L�L$hL�$H�D$pH�D$L�D$H�D$�    H��$�   �\$ H��< u~L��$�   H�5    H��   H9�|_H�|$@H9�wNL�D$8H9�u@L�D$hL�$H�D$pH�D$H�t$XH�t$H�D$`H�D$�    �\$ H�؈�$�   H��x�1����    1���Ƅ$�   ��1��m����    1��_���H��   �S���1������H��   �����1��m����    ��������������������
      z  go.string."."   �   runtime.eqstring   �  go.string.".."   �   runtime.eqstring   �  go.string."./"   �   runtime.eqstring   �  go.string."../"   �   runtime.eqstring   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   0�  "".autotmp_0820  type.bool "".autotmp_0819  type.bool "".autotmp_0818  type.string "".autotmp_0817  type.int "".autotmp_0816  type.int "".autotmp_0815  type.int "".autotmp_0814 type.string "strings.prefix·3 ?type.string strings.s·2 type.string "strings.prefix·3 _type.string strings.s·2 �type.string "".~r1  type.bool "".path  type.string  ����T� � "�
&'&�  O� Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c   :$GOROOT/src/go/build/build.go�"".ArchChar  �  �dH�%    H;a��   H��H1�H�\$`H�\$h1�H�\$pH�\$xH�    H�\$8H�D$@"   1�H�\$(H�\$0H�    H�$�    H�D$H�D$ H�l$@H�hH�l$8�=     unH�(H�D$ H�    1�H9�t)H�L$ H�    H�\$`H�D$h   H�D$pH�L$xH��H�H�    H�$H�    H�\$H�    H�\$�    H�D$�H�$H�l$�    H�D$ ��    �������
      d  \go.string."architecture letter no longer used"   �  .type.errors.errorString   �  "runtime.newobject   � (runtime.writeBarrier   �  Bgo.itab.*errors.errorString.error   �  go.string."?"   �  0type.*errors.errorString   �  type.error   �  Bgo.itab.*errors.errorString.error   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   `�  "".autotmp_0825 O0type.*errors.errorString "".autotmp_0824  0type.*errors.errorString "".~r0 ?type.error errors.text·2 type.string "".~r2 @type.error "".~r1  type.string "".goarch  type.string  ����D� � �/�  [�- Tgclocals·adb3347b296419e60da36d67f8b7ce43 Tgclocals·11d28ee4a7546638afa514476454a63e   :$GOROOT/src/go/build/build.go�"".isIdent  `  `�D$<Ar
<Zw�D$�<ar<zv�<0r<9v�<_t�<��D$��     "".~r1 type.bool "".c  type.uint8 0 0 
.+  Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�<"".(*importReader).syntaxError  �  �dH�%    H;avKH��H�D$H�h(H�� uH�-    H�h(H�-    �=     u	H�h0H���L�@0L�$H�l$�    ���    ����������������
      J  "".errSyntax   ` "".errSyntax   l (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt      "".r  *type.*"".importReader  2  p B
 
 S Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�6"".(*importReader).readByte  �  �dH�%    H;a��  H��hH�\$pH�+H�,$�    L�L$p�\$H�ވ\$GH�|$H�\$H�\$`H�|$XH�� u?I�QI�AI�IH��H��H9���   I�iH�@�3@�� uH�=    H�    H�\$`H�� t]H�-    H9�u[H�|$XH�<$H�l$`H�l$H�-    H�l$H�-    H�l$�    L�L$pH�|$X�\$ �� tH��   A�i81�@�t$xH��h�I�i(H�� u�H�|$XI�y(H�l$`�=     uI�i0��M�A0L�$H�l$�    �H�    H�$H�T$H�D$H�L$H�l$ �    L�L$pH�|$X�t$GH�T$(H�D$0H�L$8I�� tZH��H�D$HH��I�iI�IH�T$P�=     u	I�Q�����M�AL�$H�T$�    L�L$pH�|$X�t$GH�T$PH�D$H����A���    ���������
      H  0bufio.(*Reader).ReadByte   �  "".errNUL   � "".errNUL   �  io.EOF   �  io.EOF   � io.EOF   �  runtime.ifaceeq   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]uint8   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".err type.error "".c Atype.uint8 "".~r0 type.uint8 "".r  *type.*"".importReader "������ � LR1&P
	
�  #�d&`7 Tgclocals·f7309186bf9eeb0f8ece2eb16f2dc110 Tgclocals·fce3d64185acee4a98aea2303545fc5c   8$GOROOT/src/go/build/read.go�6"".(*importReader).peekByte  �
  �
dH�%    H;a��  H��@H�T$HH�j(H�� tvH�j@H��H�j@H�Z@H��'  ~TH�    H�\$0H�D$8   H�    H�$H�\$0H�\$H�D$    �    H�\$H�H�$H�KH�L$�    �D$X H��@��j H��@�� uH�$�    H�T$H�\$H��H�j(H�� u:�Z8�� u1�|$P t*��wB��	u1H�$�    H�T$H�\$H��H�j(H�� tƈJ �j @�l$XH��@À�
tʀ�t���� w��t��� t��Ҁ�/�N  H�$�    H�L$H�\$H�؀�/uL<
t-H�i(H�� u#�Y8�� uH�$�    H�L$H�\$H��<
u�H�$�    H�T$H�\$H��������*��   1҈T$/<*tbH�i(H�� u��Y8�� t)H�i(H�� uH�-    H�i(H�-    �=     u5H�i0H�$�    H�L$H�\$H���\$/H�؈T$/<*u���/�g����L�A0L�$H�l$�    H�L$H�H�i(H�� �>���H�-    H�i(H�-    �=     u	H�i0����L�A0L�$H�l$�    H�L$H�������;�R����m����    �`���(
      �  Vgo.string."go/build: import reader looping"   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  6"".(*importReader).readByte   �  6"".(*importReader).readByte   �  6"".(*importReader).readByte   �  6"".(*importReader).readByte   �  6"".(*importReader).readByte   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  6"".(*importReader).readByte   �  .runtime.writebarrierptr   �	  "".errSyntax   �	 "".errSyntax   �	 (runtime.writeBarrier   �	  .runtime.writebarrierptr   �
  0runtime.morestack_noctxt   0�  "".autotmp_0834  type.uint8 "".autotmp_0833 type.string 
"".c1 !type.uint8 "".~r1  type.uint8 "".skipSpace type.bool "".r  *type.*"".importReader (���w��
 � �|
T

@7
67
6-	3		)"-)	6]
  q<� Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·d8fdd2a55187867c76648dc792366181   8$GOROOT/src/go/build/read.go�6"".(*importReader).nextByte  �  �dH�%    H;av5H��H�\$ H�$�\$(�\$�    �\$H��H�\$ �C  �D$0H����    ������
      L  6"".(*importReader).peekByte   �  0runtime.morestack_noctxt   00  "".~r1  type.uint8 "".skipSpace type.bool "".r  *type.*"".importReader 00/ P �		 
 %+ Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�<"".(*importReader).readKeyword  �  �dH�%    H;a�U  H�� H�\$(H�$�D$�    H�t$(H�T$81�H�L$H9���   H�4$�D$ �    H�t$(H�T$8H�L$�\$H��H�\$0H9���   H��8�tBH�n(H�� uH�-    H�n(H�-    �=     u	H�n0H�� �L�F0L�$H�l$�    ��H��H�L$H9��o���H�4$�D$ �    �\$H�؀�ArV<ZwRH��   < t.H�D$(H�h(H�� uH�-    H�h(H�-    �=     u	H�h0H�� �L�@0L�$H�l$�    ��<ar<zv�<0r<9v�<_t�<�����    �    ������������������
      L  6"".(*importReader).peekByte   �  6"".(*importReader).nextByte   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  6"".(*importReader).peekByte   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0@  
"".autotmp_0839  type.uint8 "".autotmp_0836  type.int "".i type.int 
"".kw type.string "".r  *type.*"".importReader "@�?@�?@6? � H�>)*.	  %� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�8"".(*importReader).readIdent  �  �dH�%    H;a�  H��H�\$ H�$�D$�    H�L$ �\$H�؀�A��   <Z��   H��   < uBH�i(H�� uH�-    H�i(H�-    �=     u	H�i0H���L�A0L�$H�l$�    ��H�$�D$ �    H�L$ �\$H�؀�Ar<ZwH��   < t�A  ��H���<ar<zv�<0r<9v�<_t�<�����<ar<z�R���<0r<9�F���<_�>���<����;����    �������
      L  6"".(*importReader).peekByte   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  6"".(*importReader).peekByte   �  0runtime.morestack_noctxt   0  "".autotmp_0843  type.bool "".r  *type.*"".importReader 0i/0M/0E/ � <�)/*  %� Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�:"".(*importReader).readString  �  �dH�%    H�D$�H;A��  H��   H��$�   H�$�D$�    H��$�   �\$��"�8  H�XH��H�\$PH�h(H�� ��   H�$�D$ �    H��$�   �\$H�ڈ\$G��"�u  H��$�   1�H9���   H�l$PL�@L�HL9��E  L�PI)�I)�I�� tM�*H�$    L�T$xL�T$L��$�   L�D$L��$�   L�L$�    H�\$ H�\$hH�\$(H�\$pH��$�   H�H�kH�KH��H��H9�wCH�kH��H��Hk�H�H�l$pH�kH�l$h�=     uH�+H�Đ   �H�$H�l$�    ��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$�   H�� tFH��H�l$XH��H�kH�KH�T$`�=     uH��W���H�$H�T$�    H�T$`H�D$X�:������    �X8�� u)��
t$��\�;���H�$�D$ �    H��$�   � ���H�h(H�� u�H�-    H�h(H�-    �=     uH�h0�L�@0L�$H�l$�    �T$GH��$�   됀�`�  H�XH��H�\$HH�h(H�� �����H�$�D$ �    H��$�   �\$��`�u  H��$�   1�H9��~���H�l$HL�@L�HL9��E  L�PI)�I)�I�� tM�*H�$    L�T$xL�T$L��$�   L�D$L��$�   L�L$�    H�\$ H�\$hH�\$(H�\$pH��$�   H�H�kH�KH��H��H9�wCH�kH��H��Hk�H�H�l$pH�kH�l$h�=     uH�+�����H�$H�l$�    ����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$�   H�� tFH��H�l$XH��H�kH�KH�T$`�=     uH��W���H�$H�T$�    H�T$`H�D$X�:������    �X8�� �L���H�h(H�� �>���H�-    H�h(H�-    �=     u	H�h0����L�@0L�$H�l$�    H��$�   �����H�h(H�� �����H�-    H�h(H�-    �=     u	H�h0����L�@0L�$H�l$�    �u����    ����D
      b  6"".(*importReader).nextByte   �  6"".(*importReader).nextByte   �  2runtime.slicebytetostring   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  6"".(*importReader).nextByte   �	  "".errSyntax   �	 "".errSyntax   �	 (runtime.writeBarrier   �	  .runtime.writebarrierptr   �
  6"".(*importReader).nextByte   �  2runtime.slicebytetostring   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  "".errSyntax   � "".errSyntax   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".autotmp_0852  type.string "".autotmp_0851 Otype.string "".autotmp_0849  type.[]uint8 "".autotmp_0848  type.int "".autotmp_0847 /type.[]uint8 "".autotmp_0846  type.uint8 "".c �type.uint8 "".start type.int "".start �type.int "".save type.*[]string "".r  *type.*"".importReader "������
 �	 ��#	�'(�	)3	$��-:-?@?
 ( 0�T�T� Tgclocals·7e902992778eda5f91d29a3f0c115aee Tgclocals·a1435607261436f22ba8c52b7acb6d2b   8$GOROOT/src/go/build/read.go�:"".(*importReader).readImport  �  �dH�%    H;a��   H��H�\$ H�$�D$�    H�L$ �\$H�؀�.u�A  H�$H�\$(H�\$�    H��À�Ar<ZwH��   < t�H�$�    H�L$ ��<ar<zv�<0r<9v�<_t�<������    �_������������������

      L  6"".(*importReader).peekByte   �  :"".(*importReader).readString   �  8"".(*importReader).readIdent   �  0runtime.morestack_noctxt    0  "".imports type.*[]string "".r  *type.*"".importReader 0@/0?/ � 0�   %� Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/build/read.go�"".readComments  �  �dH�%    H��$H���H;A��  H��8  1�H��$P  H��$X  H��$`  1�H��$h  H��$p  H��$@  H��$H  H�\$`H�D$hH�D$xH��   H�\$p1�H9�tH�[H�-    H9��  H��   �� ��   H�XH9���   H��$�   W��    G�H��$�   H��H�� ��   W��    G�H�H�\$@H�$�D$�    H�D$@H�h(H�� u�X8�� uH�HH��L�@L9�wRH�HH�� tDH�hH��$P  H�hH��$X  H�hH��$`  H�h(H��$h  H�h0H��$p  H��8  É ��    ��V���H�T$0H��}	H�D$0   H�    H�$�    H�L$0H�D$H�D$8H�D$HH�    H�$H�L$H�L$�    H�t$H�l$ H�T$(H�L$pH�D$xH��$�   W�H����    G�H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H�L$PH��$�   H�D$XH��$   HǄ$(  ����HǄ$0  ����H�\$HH�� t,H��$�   H�\$H�l$H�-    H�,$�    H�D$8�������1�1�������    �I������������
      �  $type.*bufio.Reader   ��  runtime.duffzero   ��  runtime.duffzero   �  6"".(*importReader).peekByte   �  $runtime.panicslice   �  "type.bufio.Reader   �  "runtime.newobject   �  type.[]uint8   �  "runtime.makeslice   ��  runtime.duffzero   �
  "type.bufio.Reader   �
  (runtime.typedmemmove   �
  0runtime.morestack_noctxt   p�  "".autotmp_0868 �(type."".importReader "".autotmp_0866  $type.*bufio.Reader "".autotmp_0864  type.int "".autotmp_0863 �"type.bufio.Reader bufio.r·3 �type.io.Reader bufio.buf·2 �type.[]uint8 bufio.b·1 �$type.*bufio.Reader bufio.r·6 �$type.*bufio.Reader bufio.size·3 �type.int bufio.rd·2 �type.io.Reader bufio.rd·2 �type.io.Reader "".r �*type.*"".importReader "".~r2 Ptype.error "".~r1  type.[]uint8 "".f  type.io.Reader ""������ � ,�N�N�  �
-.�/ Tgclocals·28b6eb03a42390d78755fe1e234a72ea Tgclocals·70b96bb4883c3816d291a08b355c816f   8$GOROOT/src/go/build/read.go�"".readImports  �  �dH�%    H��$8���H;A�p  H��H  1�H��$p  H��$x  H��$�  1�H��$�  H��$�  H��$P  H��$X  H�\$`H�D$hH�D$xH��   H�\$p1�H9�tH�[H�-    H9���  H��   �� ��  H�XH9���  H��$�   W��    G�H��$�   H��H�� ��  W��    G�H�H�\$@H�$H�    H�\$H�D$   �    H�\$@H�$�    H�\$@H�$�D$�    H�D$@�\$��i��   H�$H�    H�\$H�D$   �    H�\$@H�$�D$�    H�L$@�\$��(ueH�$�D$ �    H�\$@H�$�D$�    H�L$@�\$��)t"H�i(H�� uH�$H��$h  H�\$�    �H�$�D$ �    �5���H�$H��$h  H�\$�    ����H�h(H�� uV�X8�� uMH�HH��L�@L9�w6L�HL��$p  H��$x  L��$�  1�H��$�  H��$�  H��H  ��    H�� ��   H�H(H�P0H�-    H9���   H��$�   H�$H��$�   H�T$H�-    H�l$H�-    H�l$�    H�D$@�\$ �� t?��$`   u51�H�h(H�h0H�h(H�� u!�X8�� uH�$�    H�D$@H�h(H�� t�H�� tDH�hH��$p  H�hH��$x  H�hH��$�  H�h(H��$�  H�h0H��$�  H��H  É 븉 ������x���H�T$0H��}	H�D$0   H�    H�$�    H�L$0H�D$H�D$8H�D$HH�    H�$H�L$H�L$�    H�t$H�l$ H�T$(H�L$pH�D$xH��$�   W�H����    G�H��$�   H��$�   H��$�   H��$�   H��$�   H��$   H�L$PH��$  H�D$XH��$  HǄ$8  ����HǄ$@  ����H�\$HH�� t,H��$�   H�\$H�l$H�-    H�,$�    H�D$8�3������1�1������    �k��������������<
      �  $type.*bufio.Reader   ��  runtime.duffzero   ��  runtime.duffzero   �  &go.string."package"   �  <"".(*importReader).readKeyword   �  8"".(*importReader).readIdent   �  6"".(*importReader).peekByte   �  $go.string."import"   �  <"".(*importReader).readKeyword   �  6"".(*importReader).peekByte   �  6"".(*importReader).nextByte   �  6"".(*importReader).peekByte   �  :"".(*importReader).readImport   �  6"".(*importReader).nextByte   �  :"".(*importReader).readImport   �	  $runtime.panicslice   �	  "".errSyntax   �
  "".errSyntax   �
 "".errSyntax   �
  runtime.ifaceeq   �  6"".(*importReader).readByte   �  "type.bufio.Reader   �  "runtime.newobject   �  type.[]uint8   �  "runtime.makeslice   ��  runtime.duffzero   �  "type.bufio.Reader   �  (runtime.typedmemmove   �  0runtime.morestack_noctxt   ��  ("".autotmp_0882 �type.error "".autotmp_0881 �(type."".importReader "".autotmp_0879  $type.*bufio.Reader "".autotmp_0878  type.[]uint8 "".autotmp_0877  type.int "".autotmp_0876  type.int "".autotmp_0872 �"type.bufio.Reader bufio.r·3 �type.io.Reader bufio.buf·2 �type.[]uint8 bufio.b·1 �$type.*bufio.Reader bufio.r·6 �$type.*bufio.Reader bufio.size·3 �type.int bufio.rd·2 �type.io.Reader bufio.rd·2 �type.io.Reader "".r �*type.*"".importReader "".~r4 ptype.error "".~r3 @type.[]uint8 "".imports 0type.*[]string ("".reportSyntaxError  type.bool "".f  type.io.Reader 0"��������� �	 x�N�#&",M
q


N1�D & �
�Z�.�1 Tgclocals·956d50cd930e9c0fc470cac7c8ba19b7 Tgclocals·8be1320446f57d096ee33ca6a889aca6   8$GOROOT/src/go/build/read.go�4"".(*Context).Import.func1  �  �dH�%    H��$`���H;A�}  H��   H�BH�ZH�\$XH�ZH�\$`H�Z H�+H�l$hH�kH�l$pH�� �:  H�hHH��$�   H�@PH���  H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� ��   H�$    H�\$hH�\$H�\$pH�\$H�    H�\$H�D$    H�t$XH�� txH�^@H�|$(H�H�H�KH�OH�    H�\$8H�D$@   �    H�L$HH�D$PH�\$`H��$�   H�CH��$�   �=     uH�H��   �H�$H�L$�    ���H��u�H��$�   H�,$H��$�   H�D$H�-    H�l$H�D$   �    �\$ �� t�H�t$XH�� ��  H�^@H�H�$H�KH�L$�    H�\$H��$�   H�\$H��$�   H�\$ H�\$xH�\$(H��$�   H��$�   H��H�� �`  H�5    �    HǄ$�      HǄ$�      H��H��$�   H�l$pH�kH�l$h�=     ��   H�+H��$�   H��H�� H�kH��$�   �=     ��   H�+H��$�   H��H��@H�kH�l$x�=     uvH�+H�$    H�D$H��$�   H�\$H��$�   H�\$�    H�L$ H�D$(H�\$`H��$�   H�CH��$�   �=     uH��7���H�$H�L$�    �$���H�$H�l$�    H��$�   �r���H�$H�l$�    H��$�   �3���H�$H�l$�    H��$�   ������������3���� �����    �^�����������������.
      �  go.string."gc"   �   runtime.eqstring   �  go.string."/"   �  go.string.".a"   �  *runtime.concatstring4   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  "go.string."gccgo"   �   runtime.eqstring   �  path.Split   �  """.statictmp_0886   ��  runtime.duffcopy   �	 (runtime.writeBarrier   �
 (runtime.writeBarrier   �
 (runtime.writeBarrier   �  *runtime.concatstrings   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  "runtime.morestack    �  "".autotmp_0885 �type.[]string "".autotmp_0884 �type.string "".autotmp_0883 �type.[6]string  "".pkgtargetroot �type.string "".&pkga �type.*string "".p � type.*"".Package "".elem �type.string "".dir �type.string ""������ � P�MS�CY�X 4 ��E?2�B? Tgclocals·7be4bbacbfdb05fb3044e36c22b41e8b Tgclocals·d471303acc881ec3c678ddfbe4bb4911   :$GOROOT/src/go/build/build.go�4"".(*Context).Import.func2  �  �dH�%    H;a��  H��xH��$�   H�$H��$�   H�\$H�    H�\$H�D$
   �    L��$�   �\$ �� ��  H��$�   H�|$(H�5    H�t$HH��	   L�L$0H�D$PI9��\  L��H)�L��L9��C  H)�I��H�� tM�H9��#  L�D$hL�$H�l$pH�l$H�t$H�D$�    L��$�   �\$ H��< ��   H��$�   H�|$8H�5    H�t$XH��	   L�L$@H�D$`I9���   L9���   H9���   H�|$hH�<$H�D$pH�D$H�t$H�D$�    L��$�   �\$ H��< uLI��u<H��$�   H�$L�L$H�    H�\$H�D$   �    �\$ ��$�   H��x�Ƅ$�    ��Ƅ$�   ��1���    1��H��   �1������    1������H��   ������    ���������
      f  ,go.string."/testdata/"   �   strings.Contains   �  *go.string."/testdata"   �   runtime.eqstring   �  *go.string."testdata/"   �   runtime.eqstring   �  (go.string."testdata"   �   runtime.eqstring   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   0�  "".autotmp_0902  type.bool "".autotmp_0900  type.string "".autotmp_0899  type.int "".autotmp_0898  type.int "".autotmp_0897  type.int "".autotmp_0896 type.string "strings.prefix·3 ?type.string strings.s·2 type.string "strings.suffix·3 _type.string strings.s·2 �type.string "".~r1  type.bool "".sub  type.string  ����M� � ��  E� Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c   :$GOROOT/src/go/build/build.go�4"".(*Context).Import.func3  �$  �$dH�%    H��$����H;A��  H��  H�rH�ZH�H�CH�Z H�+H��$  H�kH��$  H�Z0H�\$PH�Z8H�\$HH�Z@H�\$hH�t$XH�4$H��$�  H�\$H��$�  H�\$H��$�   H�L$H��$�   H�D$ �    L�T$(L�L$0�\$8�� �  L��$�   L��$�   L��$�   H�=    H��$   H��   L��$�   H��$  I9���  L9���  H9���  L��$0  L�$H��$8  H�D$H�|$H�D$�    L��$�   L��$�   �\$ H��< �k  L�$L�L$H�    H�\$H�D$
   �    �\$ �� �:  H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hH�-    H�h H�-    H�h(HǄ$H     HǄ$P     H��$@  H��$�  H�hH��$�  �=     ��  H�(H��$�   H��H��H�kH��$�   �=     �B  H�+H�\$XH�$H�D$H��$H  H�\$H��$P  H�\$�    H�L$ H�D$(H�\$XH�$H��$�   H�L$H��$�   H�D$�    �\$�� ��  H�    H�$�    H�D$H�� ��  HǄ$H     HǄ$P     H��$@  H��$�   H�hH��$�   �=     �K  H�(H��$  H��H��H�kH��$  �=     �  H�+H�\$XH�$H�D$H��$H  H�\$H��$P  H�\$�    H�L$ H�D$(H�\$XH�$H��$   H�L$H��$(  H�D$�    �\$�� �H  H�\$XH�$H��$   H�\$H��$(  H�\$�    �\$�� �  H�\$PH��$(  H�kH��$   �=     ��  H�+H��$X  H��H�-    H�+H�-    H�kH�-    H�kH�-    H�kH�-    H�k H�-    H�k(HǄ$H     HǄ$P     H��$@  H��$�   H�kH��$�   �=     �.  H�+H��$  H��H�� H�kH��$  �=     ��  H�+H�$H��$H  H�\$H��$P  H�\$�    H�T$H�t$ L�    I��   1�H�\$pH�\$xH��$�   H��$�   H��$�   L��$�   L��$�   L��$�   H��$�   L��$�   L9��N  I9��>  M9��.  H��$0  H�$L��$8  L�T$L�D$L�T$�    L��$�   H��$�   H��$�   �\$ H��< ��   H��I9���   L)�I��H�� tO�L��H��H�\$PH�� ��   H�D$xH�CHH�T$p�=     ulH�S@H�\$P��$�  @���   H�\$PH��$�  H�kXH��$�  �=     uH�kPH�T$HH���Ƅ$�  H�Ĉ  �L�CPL�$H�l$�    ��L�C@L�$H�T$�    넉�b����    H���D���1������    1�����H�$H�l$�    H��$@  � ���H�$H�l$�    H��$@  ����H�$H�l$�    ����H�\$hH�H�CH�KH��H��H9���   H�kH��H��Hk�H�H��$(  H�kH��$   �=     urH�+H��$�   H�$H��$�   H�\$H�    H�\$H�D$   �    H�D$ H�� }Ƅ$�   H�Ĉ  �H��$�   H9�wH��$�   ������    H�$H�l$�    �H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�D$0H�L$8H�\$hH��H�D$@H��H�kH�KH�T$`�=     uH������H�$H�T$�    H�T$`H�D$@�����H�$H�l$�    H��$@  �����H�$H�l$�    H��$@  ����� �R��������H�$H�l$�    H��$@  ����H�$H�l$�    H��$@  �`���Ƅ$�   H�Ĉ  �1��v����    1��h����    ��������|
      �  ."".(*Context).hasSubdir   �   go.string."src/"   �   runtime.eqstring   �  ,go.string."/testdata/"   �   strings.Contains   �  type.[3]string   �  "runtime.newobject   �  """.statictmp_0922   � """.statictmp_0922   �  """.statictmp_0922   �0 """.statictmp_0922   �@ """.statictmp_0922   �P """.statictmp_0922   � (runtime.writeBarrier   �	 (runtime.writeBarrier   �
  ,"".(*Context).joinPath   �
  &"".(*Context).isDir   �  type.[2]string   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   �  ,"".(*Context).joinPath   �  &"".(*Context).isDir   �  "".hasGoFiles   � (runtime.writeBarrier   �  """.statictmp_0927   � """.statictmp_0927   �  """.statictmp_0927   �0 """.statictmp_0927   �@ """.statictmp_0927   �P """.statictmp_0927   � (runtime.writeBarrier   � (runtime.writeBarrier   �  path.Join   �   go.string."src/"   �   runtime.eqstring   � (runtime.writeBarrier   � (runtime.writeBarrier   �       �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   � (runtime.writeBarrier   �  go.string."/"   �  "strings.LastIndex   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  (runtime.writeBarrier   �!  .runtime.writebarrierptr   �!  .runtime.writebarrierptr   �!  .runtime.writebarrierptr   �"  .runtime.writebarrierptr   �"  .runtime.writebarrierptr   �#  $runtime.panicslice   �#  "runtime.morestack   @�  B"".autotmp_0929 _type.[3]string "".autotmp_0928  type.*[3]string "".autotmp_0926  type.[]string "".autotmp_0924  type.[]string "".autotmp_0921 �type.[]string "".autotmp_0918  type.int "".autotmp_0917  type.string "".autotmp_0916  type.int "".autotmp_0915  type.int "".autotmp_0914  type.int "".autotmp_0913  type.string "".autotmp_0910  type.bool "".autotmp_0909  type.bool "".autotmp_0908 �type.string "".&tried ��type.*struct { vendor []string; goroot string; gopath []string } "".setPkga �type.func() "".p � type.*"".Package "".path �type.string "".srcDir �type.string "".ctxt � type.*"".Context "strings.prefix·3 �type.string strings.s·2 �type.string "".~r0 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "".dir �type.string "".vendor �type.string "".sub �type.string "".~r2 0type.bool "".isGoroot  type.bool "".root  type.string <"����������� � ��	gQ��6�l)�&
aP8
!"~=6 l ����2���-�:&K� Tgclocals·75ee4963a64d57666eac9d22b87e7339 Tgclocals·68281ae9cb2c0df5f0c33d324dd29c1b   :$GOROOT/src/go/build/build.go�4"".(*Context).Import.func4  �  �dH�%    H;a�e  H��hH�BH�ZH�\$HH�ZH�+H�l$XH�kH�l$`H�(H�� uH�l$pH�(H�l$x�=     �  H�hH�\$HH��(  H��0  H��8  H��H��H9�wCH��0  H��H��Hk�H�H�l$`H�kH�l$X�=     uH�+H��h�H�$H�l$�    ��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�D$0H�L$8H�\$HH�� tWH��H�D$@H��H��0  H��8  H�T$P�=     uH��(  �S���L��(  L�$H�T$�    H�T$PH�D$@�/�����L�@L�$H�l$�    ������    �~�����������������
      � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  "runtime.morestack    �  "".name type.string "".p ? type.*"".Package "".err  type.error "������ � 2�
9	S�  �&b%" Tgclocals·7e902992778eda5f91d29a3f0c115aee Tgclocals·66499ec09befdf27c68e3e35878ba2c7   :$GOROOT/src/go/build/build.go�"".init  �  �dH�%    H��$����H;A�&  H���  �    �� t�    ��uH���  ��    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     �E  H�    1�H��}gH�    H�$H�    H�\$H�    H��Hk�H�H�\$H�    H��H��$�   Hk�H�H�\$H�D$�    H��$�   H��H��|��    H��$   H���    H��$   H�-    H�l$H�\$H�    H�$�    H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     �:  H�    H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     ��  H�    �    H�$H��$�   H�\$H��$�   H�    H�$�    H�D$H�-    H�(H�-    H�hH�-    H�hH�-    H�hHǄ$�      HǄ$�      H��$�   H��$�   H�hH��$�   �=     �  H�(H�$H��$�   H�\$H��$�   H�\$�    H�\$ H�    H�\$�=     ��   H�    H�    H�$H�D$   �    H�\$H�    H�\$�=     ulH�    H�    H�$H�D$   �    H�\$H�    H�\$�=     uH�    �    �    H���  �H�-    H�,$H�\$�    ��H�-    H�,$H�\$�    �H�-    H�,$H�\$�    �0���H�$H�l$�    H��$�   �����H�-    H�,$H�\$�    ����H�-    H�,$H�\$�    ����H�-    H�,$H�\$�    �����    ��������̤
      J  "".initdone·   b  "".initdone·   �  "runtime.throwinit   � "".initdone·   �  bytes.init   �  fmt.init   �  go/ast.init   �  go/doc.init   �  go/parser.init   �  go/token.init   �  io.init   �  io/ioutil.init   �  log.init   �  os.init   �  path.init   �  $path/filepath.init   �  runtime.init   �  strconv.init   �  strings.init   �  unicode.init   �  bufio.init   �  (type.map[string]bool   �  runtime.makemap   � (runtime.writeBarrier   �  "".cgoEnabled   �  (type.map[string]bool   �  "".cgoEnabled   �  """.statictmp_0939   �  """.statictmp_0939   �  $runtime.mapassign1   �  """.defaultContext   ��  runtime.duffcopy   �  "".Default   �  type."".Context   �  (runtime.typedmemmove   �  (type.map[string]bool   �  runtime.makemap   � (runtime.writeBarrier   �  "".knownOS   �  (type.map[string]bool   �  runtime.makemap   � (runtime.writeBarrier   �  "".knownArch   �  runtime.GOROOT   �  type.[2]string   �	  "runtime.newobject   �	  """.statictmp_0942   �	 """.statictmp_0942   �	  """.statictmp_0942   �	0 """.statictmp_0942   �
 (runtime.writeBarrier   �  $path/filepath.Join   � "".ToolDir   � (runtime.writeBarrier   �  "".ToolDir   �  0go.string."syntax error"   �  errors.New   �  "".errSyntax   � (runtime.writeBarrier   � "".errSyntax   �  Fgo.string."unexpected NUL in input"   �  errors.New   �  "".errNUL   � (runtime.writeBarrier   � "".errNUL   �  "".init.1   � "".initdone·   � "".errNUL   �  .runtime.writebarrierptr   � "".errSyntax   �  .runtime.writebarrierptr   �  "".ToolDir   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  "".knownArch   �  .runtime.writebarrierptr   �  "".knownOS   �  .runtime.writebarrierptr   �  "".cgoEnabled   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".autotmp_0941 �type.[]string "".autotmp_0940 �type.int "".autotmp_0938 �type.string "".autotmp_0937 �type."".Context ."�������� 2��ti v��Do5>�DD��::'('&�����   B���"M Tgclocals·7d2d5fca80364273fb07d5820a76fef4 Tgclocals·826f148c2b9ed682d2ed28d3c55a6368   >$GOROOT/src/go/build/syslist.go:$GOROOT/src/go/build/build.go8$GOROOT/src/go/build/read.go�(type..hash.[8]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0948 type.int "".autotmp_0947 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[8]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�$type..eq.[8]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_0952 ?type.string "".autotmp_0951 type.string "".autotmp_0950 _type.int "".autotmp_0949 Otype.int "".~r2  type.bool "".q type.*[8]string "".p  type.*[8]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�(type..hash.[2]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0954 type.int "".autotmp_0953 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[2]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�$type..eq.[2]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_0958 ?type.string "".autotmp_0957 type.string "".autotmp_0956 _type.int "".autotmp_0955 Otype.int "".~r2  type.bool "".q type.*[2]string "".p  type.*[2]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�(type..hash.[6]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0960 type.int "".autotmp_0959 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[6]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�$type..eq.[6]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_0964 ?type.string "".autotmp_0963 type.string "".autotmp_0962 _type.int "".autotmp_0961 Otype.int "".~r2  type.bool "".q type.*[6]string "".p  type.*[6]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�4type..hash.[5]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0966 type.int "".autotmp_0965 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[5]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�0type..eq.[5]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0970 ?"type.interface {} "".autotmp_0969 "type.interface {} "".autotmp_0968 _type.int "".autotmp_0967 Otype.int "".~r2  type.bool "".q *type.*[5]interface {} "".p  *type.*[5]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�(type..hash.[3]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0972 type.int "".autotmp_0971 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[3]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�$type..eq.[3]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_0976 ?type.string "".autotmp_0975 type.string "".autotmp_0974 _type.int "".autotmp_0973 Otype.int "".~r2  type.bool "".q type.*[3]string "".p  type.*[3]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�4type..hash.[1]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0978 type.int "".autotmp_0977 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[1]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�0type..eq.[1]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0982 ?"type.interface {} "".autotmp_0981 "type.interface {} "".autotmp_0980 _type.int "".autotmp_0979 Otype.int "".~r2  type.bool "".q *type.*[1]interface {} "".p  *type.*[1]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�4type..hash.[2]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0984 type.int "".autotmp_0983 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[2]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�0type..eq.[2]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0988 ?"type.interface {} "".autotmp_0987 "type.interface {} "".autotmp_0986 _type.int "".autotmp_0985 Otype.int "".~r2  type.bool "".q *type.*[2]interface {} "".p  *type.*[2]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go��type..hash.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } �  �dH�%    H;avvH�� H�\$(H�$H�<$ tYH�\$0H�\$H�D$    �    H�D$H�\$(H�$H�<$ t#H�$ H�D$0H�D$�    H�\$H�\$8H�� É%    �ԉ%    ��    �q����
      n  runtime.memhash   �  runtime.strhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  �type.*struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } @_?@? � � 
 6Z Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go��type..eq.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } �  �dH�%    H;a��   H��HH�\$PH�$H�<$ ��   H�\$XH�\$H�|$ ��   H�D$    �    �\$�� u
�D$` H��H�H�\$PH�� tnH�s H�K(H�\$XH�� tWH�S H�C(H9�u@H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� t
�D$`H��H��D$` H��HÉ륉뎉%    �U����%    �3����    �������������������
      �   runtime.memequal   �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  
"".autotmp_0991 ?type.string "".autotmp_0990 type.string "".~r2  type.bool "".q �type.*struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } "".p  �type.*struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } 6�K��j��	�� � � �  J� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go��type..hash.struct { F uintptr; badGoError *error; p *"".Package; name string } �  �dH�%    H;avvH�� H�\$(H�$H�<$ tYH�\$0H�\$H�D$   �    H�D$H�\$(H�$H�<$ t#H�$H�D$0H�D$�    H�\$H�\$8H�� É%    �ԉ%    ��    �q����
      n  runtime.memhash   �  runtime.strhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  �type.*struct { F uintptr; badGoError *error; p *"".Package; name string } @_?@? � � 
 6Z Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go��type..eq.struct { F uintptr; badGoError *error; p *"".Package; name string } �  �dH�%    H;a��   H��HH�\$PH�$H�<$ ��   H�\$XH�\$H�|$ ��   H�D$   �    �\$�� u
�D$` H��H�H�\$PH�� tnH�sH�K H�\$XH�� tWH�SH�C H9�u@H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� t
�D$`H��H��D$` H��HÉ륉뎉%    �U����%    �3����    �������������������
      �   runtime.memequal   �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  
"".autotmp_0994 ?type.string "".autotmp_0993 type.string "".~r2  type.bool "".q �type.*struct { F uintptr; badGoError *error; p *"".Package; name string } "".p  �type.*struct { F uintptr; badGoError *error; p *"".Package; name string } 6�K��j��	�� � � �  J� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�Ltype..hash.struct { a string; b bool } �  �dH�%    H;avvH�� H�\$(H�$H�<$ tYH�\$0H�\$�    H�D$H�\$(H�$H�<$ t,H�$H�D$0H�D$H�D$   �    H�\$H�\$8H�� É%    �ˉ%    ��    �q����
      \  runtime.strhash   �  runtime.memhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  Btype.*struct { a string; b bool } @_?@? � � 
 -c Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�Htype..eq.struct { a string; b bool } �  �dH�%    H;a��   H��HH�\$PH�� ��   H�3H�KH�\$XH�� txH�H�CH9�ubH�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� t,H�l$P�]L�D$XA�h@8�t
�D$` H��H��D$`H��H��D$` H��HÉ넉�k����    �;��������������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  
"".autotmp_0996 ?type.string "".autotmp_0995 type.string "".~r2  type.bool "".q Btype.*struct { a string; b bool } "".p  Btype.*struct { a string; b bool } 8����	��	��� � � 
 ke Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/build/build.go�Ttype..hash.[24]struct { a string; b bool } �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��Hk�H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  Ltype..hash.struct { a string; b bool }   �  0runtime.morestack_noctxt   0P  
"".autotmp_0998 type.int "".autotmp_0997 type.int "".~r2  type.uintptr "".h type.uintptr "".p  Jtype.*[24]struct { a string; b bool } PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/build/build.go�Ptype..eq.[24]struct { a string; b bool } �  �dH�%    H;a�  H��h1�H�D$(   H�l$(H9���   H�D$0H�L$pH�� ��   H�\$xH��Hk�H�H�� ��   H��Hk�H�H�L$@H�� ��   H�1H�IH�\$8H�� ��   H�H�CH9�uqH�t$XH�4$H�L$`H�L$H�T$HH�T$H�D$PH�D$�    �\$ �� t;H�l$@�]L�D$8A�h@8�u#H�D$0H��H�l$(H9��4���Ƅ$�   H��h�Ƅ$�    H��hÉ�o�����R�����2���������    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1004 ?type.string "".autotmp_1003 type.string "".autotmp_1002 _Btype.*struct { a string; b bool } "".autotmp_1001 OBtype.*struct { a string; b bool } "".autotmp_1000 type.int "".autotmp_0999 otype.int "".~r2  type.bool "".q Jtype.*[24]struct { a string; b bool } "".p  Jtype.*[24]struct { a string; b bool } ,������� � �  �� Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·34eab47d33fa46b254c22cdccfd2dc77   :$GOROOT/src/go/build/build.go�Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·d98f60bd8519d0c68364b2a1d83af357             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·d98f60bd8519d0c68364b2a1d83af357             �"go.string.hdr."/"                       go.string."/"   �go.string."/"   /  �Tgclocals·895d0569a38a56443b84805daa09d838              �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �Tgclocals·b4e92317a1ad7fa1f283390980fe4780 (  (                 �Tgclocals·dd9ae044070cfdff36caf84fd74b60b9 (  (                �Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c      
        �Tgclocals·12ab5efd4c34ee1072eaafe77351d565             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·6d46c0650eba7dbebc0db316e0e0cf3b             �><go.itab.*os.File.io.ReadCloser     �Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60                   �Tgclocals·5cbd57cf8f9b35eac9551b20a42afe1f                  �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �"go.string.hdr."~"                       go.string."~"   �go.string."~"   ~  �Tgclocals·e2234b98cb6fbb40cb1b6c335fab0a3e 8  8           �  !�  !   �   �Tgclocals·087344e727b14a841dc6a2833d52f059 8  8                      �&go.string.hdr."src"                       go.string."src"   �go.string."src"   src  �Tgclocals·605a1b837cd4aeeb8235060aa13f27b7 `  `
                           	  	    �Tgclocals·cffcb3fa139580cffca8ac28af4ff263 `  `
                                     �,go.string.hdr."GOARCH"                       $go.string."GOARCH"   �$go.string."GOARCH"   GOARCH  �*go.string.hdr."amd64"                       "go.string."amd64"   �"go.string."amd64"   amd64  �(go.string.hdr."GOOS"                        go.string."GOOS"   � go.string."GOOS"   
GOOS  �*go.string.hdr."linux"                       "go.string."linux"   �"go.string."linux"   linux  �,go.string.hdr."GOPATH"                       $go.string."GOPATH"   �$go.string."GOPATH"   GOPATH  �$go.string.hdr."gc"                       go.string."gc"   �go.string."gc"   gc  �*go.string.hdr."go1.1"                       "go.string."go1.1"   �"go.string."go1.1"   go1.1  �*go.string.hdr."go1.2"                       "go.string."go1.2"   �"go.string."go1.2"   go1.2  �*go.string.hdr."go1.3"                       "go.string."go1.3"   �"go.string."go1.3"   go1.3  �*go.string.hdr."go1.4"                       "go.string."go1.4"   �"go.string."go1.4"   go1.4  �*go.string.hdr."go1.5"                       "go.string."go1.5"   �"go.string."go1.5"   go1.5  �*go.string.hdr."go1.6"                       "go.string."go1.6"   �"go.string."go1.6"   go1.6  �6go.string.hdr."CGO_ENABLED"                       .go.string."CGO_ENABLED"   �.go.string."CGO_ENABLED"    CGO_ENABLED  �"go.string.hdr."0"                       go.string."0"   �go.string."0"   0  �"go.string.hdr."1"                       go.string."1"   �go.string."1"   1  �Tgclocals·b747f90b0df18c3781c6f6b1a3b90488 @  @   !           �*%�   �*%�    �Tgclocals·7353ec067a80b85e773ae30131808ed8 (  (                   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·b4c25e9b09fd0cf9bb429dcefe91c353             �(go.string.hdr."main"                        go.string."main"   � go.string."main"   
main  �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �"go.string.hdr."."                       go.string."."   �go.string."."   .  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·b60dc0a6046c556b02baa766a3fd5a27             �`go.string.hdr."no buildable Go source files in "                        Xgo.string."no buildable Go source files in "   �Xgo.string."no buildable Go source files in " P  Bno buildable Go source files in   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �pgo.string.hdr."found packages %s (%s) and %s (%s) in %s"             (          hgo.string."found packages %s (%s) and %s (%s) in %s"   �hgo.string."found packages %s (%s) and %s (%s) in %s" `  Rfound packages %s (%s) and %s (%s) in %s  �Tgclocals·345f1bd1394e1f5bdb891635a73ee227 (  (           �  �  �Tgclocals·cb395d89503762333b1bfb09ba74eb12 (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �>Lgo.itab.*"".MultiplePackageError.error     �>6go.itab.*"".NoGoError.error     �\go.string.hdr."import %q: invalid import path"                       Tgo.string."import %q: invalid import path"   �Tgo.string."import %q: invalid import path" @  >import %q: invalid import path  �"go.string.hdr."_"                       go.string."_"   �go.string."_"   _  �*go.string.hdr."gccgo"                       "go.string."gccgo"   �"go.string."gccgo"   gccgo  �4go.string.hdr."pkg/gccgo_"             
          ,go.string."pkg/gccgo_"   �,go.string."pkg/gccgo_"    pkg/gccgo_  �(go.string.hdr."pkg/"                        go.string."pkg/"   � go.string."pkg/"   
pkg/  �\go.string.hdr."import %q: unknown compiler %q"                       Tgo.string."import %q: unknown compiler %q"   �Tgo.string."import %q: unknown compiler %q" @  >import %q: unknown compiler %q  �$go.string.hdr.".."                       go.string.".."   �go.string.".."   ..  �$go.string.hdr."./"                       go.string."./"   �go.string."./"   ./  �&go.string.hdr."../"                       go.string."../"   �go.string."../"   ../  �~go.string.hdr."import %q: import relative to unknown directory"             /          vgo.string."import %q: import relative to unknown directory"   �vgo.string."import %q: import relative to unknown directory" `  `import %q: import relative to unknown directory  �lgo.string.hdr."import %q: cannot import absolute path"             &          dgo.string."import %q: cannot import absolute path"   �dgo.string."import %q: cannot import absolute path" P  Nimport %q: cannot import absolute path  �Dgo.string.hdr."\t%s (vendor tree)"                       <go.string."\t%s (vendor tree)"   �<go.string."\t%s (vendor tree)" 0  $	%s (vendor tree)  �(go.string.hdr."\t%s"                        go.string."\t%s"   � go.string."\t%s"   	%s  �Fgo.string.hdr."\t%s (from $GOROOT)"                       >go.string."\t%s (from $GOROOT)"   �>go.string."\t%s (from $GOROOT)" 0  &	%s (from $GOROOT)  �Fgo.string.hdr."\t($GOROOT not set)"                       >go.string."\t($GOROOT not set)"   �>go.string."\t($GOROOT not set)" 0  &	($GOROOT not set)  �Fgo.string.hdr."\t%s (from $GOPATH)"                       >go.string."\t%s (from $GOPATH)"   �>go.string."\t%s (from $GOPATH)" 0  &	%s (from $GOPATH)  �Fgo.string.hdr."\t($GOPATH not set)"                       >go.string."\t($GOPATH not set)"   �>go.string."\t($GOPATH not set)" 0  &	($GOPATH not set)  �$go.string.hdr."\n"                       go.string."\n"   �go.string."\n"   
  �jgo.string.hdr."cannot find package %q in any of:\n%s"             $          bgo.string."cannot find package %q in any of:\n%s"   �bgo.string."cannot find package %q in any of:\n%s" P  Jcannot find package %q in any of:
%s  �&go.string.hdr."pkg"                       go.string."pkg"   �go.string."pkg"   pkg  �&go.string.hdr."bin"                       go.string."bin"   �go.string."bin"   bin  �&go.string.hdr.".go"                       go.string.".go"   �go.string.".go"   .go  �&go.string.hdr.".hh"                       go.string.".hh"   �go.string.".hh"   .hh  �$go.string.hdr.".h"                       go.string.".h"   �go.string.".h"   .h  �$go.string.hdr.".S"                       go.string.".S"   �go.string.".S"   .S  �$go.string.hdr.".c"                       go.string.".c"   �go.string.".c"   .c  �$go.string.hdr.".s"                       go.string.".s"   �go.string.".s"   .s  �$go.string.hdr.".m"                       go.string.".m"   �go.string.".m"   .m  �&go.string.hdr.".cc"                       go.string.".cc"   �go.string.".cc"   .cc  �(go.string.hdr.".hpp"                        go.string.".hpp"   � go.string.".hpp"   
.hpp  �(go.string.hdr.".cpp"                        go.string.".cpp"   � go.string.".cpp"   
.cpp  �(go.string.hdr.".cxx"                        go.string.".cxx"   � go.string.".cxx"   
.cxx  �*go.string.hdr.".swig"                       "go.string.".swig"   �"go.string.".swig"   .swig  �(go.string.hdr.".hxx"                        go.string.".hxx"   � go.string.".hxx"   
.hxx  �*go.string.hdr.".syso"                       "go.string.".syso"   �"go.string.".syso"   .syso  �0go.string.hdr.".swigcxx"                       (go.string.".swigcxx"   �(go.string.".swigcxx"    .swigcxx  �:go.string.hdr."documentation"                       2go.string."documentation"   �2go.string."documentation"    documentation  �0go.string.hdr."_test.go"                       (go.string."_test.go"   �(go.string."_test.go"    _test.go  �*go.string.hdr."_test"                       "go.string."_test"   �"go.string."_test"   _test  �dgo.string.hdr."%s:%d: cannot parse import comment"             "          \go.string."%s:%d: cannot parse import comment"   �\go.string."%s:%d: cannot parse import comment" P  F%s:%d: cannot parse import comment  �~go.string.hdr."found import comments %q (%s) and %q (%s) in %s"             /          vgo.string."found import comments %q (%s) and %q (%s) in %s"   �vgo.string."found import comments %q (%s) and %q (%s) in %s" `  `found import comments %q (%s) and %q (%s) in %s  �~go.string.hdr."%s: parser returned invalid quoted string: <%s>"             /          vgo.string."%s: parser returned invalid quoted string: <%s>"   �vgo.string."%s: parser returned invalid quoted string: <%s>" `  `%s: parser returned invalid quoted string: <%s>  �"go.string.hdr."C"                       go.string."C"   �go.string."C"   C  �fgo.string.hdr."use of cgo in test %s not supported"             #          ^go.string."use of cgo in test %s not supported"   �^go.string."use of cgo in test %s not supported" P  Huse of cgo in test %s not supported  �&go.string.hdr."cgo"                       go.string."cgo"   �go.string."cgo"   cgo  �Tgclocals·5391224ff1aeba9fa698864a89676656 �F  �Fq   :                                                            �a       ��;  )��                     �a       ��;  )��                     �a     ��;  )��                     �a      ��;  )��             �       �a       ��;  )��            �       �c       ��;  )��             �       �a       ��;  )��            �       �a       ��;  )��             �       �a     ��;  )��             �       �a      ��;  )��             �       �a       ��; x)��             �       �a       ��; x)��              �       �a       ��; x)��             �       �a     ��; x)��             �       �a      ��; x)��             �       �a       ��; x)��             �       �a       ��; x)��             �       �a       ��; x)��             �       �a       ��; x)��            �       �a       ��; x)��            �       �a       ��; x)��            �       �a      ��; x)��            �       �a       ��; x)��             �       �a       ��; x)��             �       �a      ��; x)��             �      �a       ��; x)��            �       �a       ��; x)��            �       �a  �    ��; x)��            �       �a       ��; x)��            �    �  �a       ��; x)��             �       �a       ��; x)��     @       �       �a @     ��; x)��     @      �       �a @     ��; x)��             �       �a @     ��; x)��             �       �a @     ��; x)��             �      �a @     ��; x)��             �      �a @    ��; x)��          � �       �a       ��; x)��          � �       �a       ��; x)��          � �      �a       ��; x)��          � �      �a       ��; x)��            �      �a       ��; x)��            �       �a       ��; x)��           � �       �a       ��; x)��             �       �a       ��; x)��             �       �a       ��; x)��             � (    �a      ��; x)��             � (    �a      ��; x)��            � (    �a      ��; x)��    �       � (    �a      ��;�z)�� UU�      � (    �a      ��;�z)�� UU�     � (   ��a       ��;�z)�� UU�     � (    �a       ��;�z)�� UU�     ��(    �a       ��;�z)�� UU�M     ��(   �a       ��;�z)�� UU��     ��(    �a       ��;�z)�� UU�M     ���    �c      ��;�z)�� UU�M     ���    �a      ��;�z)�� UU�     ��(    �a       ��;�z)�� UU�M     ���    �a    � ��;�z)�� UU��M     ���    �a      ��;�z)�� UU          �      �a       ��;�z)�� UU��M     ���    �a      ��;�z)�� UU��M@    ���    �a      ��;�z)�� UU��M@    ���    �a      ��;�z)�� UU��M@    ���    �a      ��;�z)�� UU��M@    ���    �a      ��;�z)�� UU��M     ���    �a      ��;�z)�� UU���     ���    �a      ��;�z)�� UU��M     ���    �a       ��;�z)�� UU��M     ���    �a      ��;�z)�� UU��M     ���    �a       ��;�z)�� UU��M     ���    �a       ��;�z)�� UU��M     ���    �a       ��;�z)�� UU��M     ���    ��     ��;�z)�� UU��M     ���    ��      ��;�z)�� UU�]   ���    �a       ��;�z)�� UU�]    ���    ��      ��;�z)�� UU�]    ���    ��       ��;�z)�� UU�]    ���    ��       ��;�z)�� UU�]    ���    ��    @  ��;�z)�� UU�]    ���    ��       ����z)�� UU�]    ���    ��      ��;�z)�� UU�]    ���    �a       ��;�z)�� UU�]    ���    ��      ��;�z)�� UU�]    ���    ��       ��;�z)�� UU�]    ���    �a       ��;�z)�� UU�     ��(    ��       ��;�z)�� UU         �      �a       ��;�z)�� UU        �      �a       ��;�z)�� UU�       �      �a       ��;�z)���UU�      �      �a       ��;�z)���UU��      �      �a       ��;�z)���UU�       �      �a       ��;�z)�� UU�       �      �a       ��;�z)�� UU�      �      �a       ��;�z)�� UU�        �      �a       ��;�z)�� UU�       �      �a       ��;�z)�� UU         �      �a       ��;�z)�� UU        �      �a       ��;�z)�� UU         �      �a      ��;�z)�� UU         �      �a   $   ��;�z)�� UU         �      �a       ��;�z)�� UU        �      �a 
    ��; x)��            �       �a 
     ��; x)��            �       �c      ��; x)��             �       �a     ��; x)��             �       �a      ��; x)��             �       �c       ��; x)��             �       �a       ��; x)��             �       �a     ��; x)��             �       �a      ��; x)��     �Tgclocals·3b32eac464325adfcb2e0feeafb27ba3 �  �q   	                                                                                                                                                                                                                                                                                                                                                       �Tgclocals·80ce1eebd7f944e81966bdd86878cedc (  (          a       �Tgclocals·14c16763214c88f6ebc22b4b638329b7 (  (                �.go.string.hdr."package"                       &go.string."package"   �&go.string."package"   package  �,go.string.hdr."import"                       $go.string."import"   �$go.string."import"   import  �Tgclocals·423fcdc350b935457e47f75dd5e63926 (  (                  �Tgclocals·adb3347b296419e60da36d67f8b7ce43 (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a             �Tgclocals·69c1753bd5f81501d95132d08af04464           �Tgclocals·b4015c155c4a804136b8d2d3fde81a78        	      A    �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·a043b57aa077fd78befe739904a3c363             �6go.string.hdr."read %s: %v"                       .go.string."read %s: %v"   �.go.string."read %s: %v"    read %s: %v  �Tgclocals·8464a0493338a790ce587fd837b5331f h  h                @                 0    D�  D�  � �Tgclocals·d644b00c61b0153799eb59e0efc3a880 h  h      K   Ki  Ki  Ki  K  K  K	  K  Ki  K	  K	   �Tgclocals·8744fb04fbd6f74dba2601338d86fe97 0  0          �  �      �Tgclocals·9f4747e6338c5bdd4db417363b8a0d83 0  0                   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5998daf4e6d23f69cd931cd9519af48e             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a             �,go.string.hdr."+build"                       $go.string."+build"   �$go.string."+build"   +build  �Tgclocals·6c1e86c4f55eb0f4f23b9aeed94efe32 @  @                     @  !    �Tgclocals·689482aa6db86c01fa54c72fbbe58e52 @  @                         �(go.string.hdr."#cgo"                        go.string."#cgo"   � go.string."#cgo"   
#cgo  �"go.string.hdr.":"                       go.string.":"   �go.string.":"   :  �Rgo.string.hdr."%s: invalid #cgo line: %s"                       Jgo.string."%s: invalid #cgo line: %s"   �Jgo.string."%s: invalid #cgo line: %s" @  4%s: invalid #cgo line: %s  �^go.string.hdr."%s: malformed #cgo argument: %s"                       Vgo.string."%s: malformed #cgo argument: %s"   �Vgo.string."%s: malformed #cgo argument: %s" @  @%s: malformed #cgo argument: %s  �.go.string.hdr."LDFLAGS"                       &go.string."LDFLAGS"   �&go.string."LDFLAGS"   LDFLAGS  �,go.string.hdr."CFLAGS"                       $go.string."CFLAGS"   �$go.string."CFLAGS"   CFLAGS  �0go.string.hdr."CPPFLAGS"                       (go.string."CPPFLAGS"   �(go.string."CPPFLAGS"    CPPFLAGS  �0go.string.hdr."CXXFLAGS"                       (go.string."CXXFLAGS"   �(go.string."CXXFLAGS"    CXXFLAGS  �4go.string.hdr."pkg-config"             
          ,go.string."pkg-config"   �,go.string."pkg-config"    pkg-config  �Rgo.string.hdr."%s: invalid #cgo verb: %s"                       Jgo.string."%s: invalid #cgo verb: %s"   �Jgo.string."%s: invalid #cgo verb: %s" @  4%s: invalid #cgo verb: %s  �Tgclocals·456125ec998d6bb6d5850305cab89579 �  �   :           B       B        P � �  P   �B      G      F       G      B                          B       �Tgclocals·5f7cd344685fbb4cd325c2c2d65d66f9 �  �                                                    �2go.string.hdr."${SRCDIR}"             	          *go.string."${SRCDIR}"   �*go.string."${SRCDIR}"    ${SRCDIR}  �Tgclocals·6347b58243cc1c5f8f735d259ec00f70 (  (          !        �Tgclocals·776d9d553b2634d9ea530b3c76543df4 (  (                �Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60                   �Tgclocals·f47057354ec566066f8688a4970cff5a                  �>Bgo.itab.*errors.errorString.error     �<go.string.hdr."unclosed quote"                       4go.string."unclosed quote"   �4go.string."unclosed quote"    unclosed quote  �Fgo.string.hdr."unfinished escaping"                       >go.string."unfinished escaping"   �>go.string."unfinished escaping" 0  (unfinished escaping  �Tgclocals·3766546ec9671d5836402e8fa0c9f6e2 P  P              	  
    �        �Tgclocals·80238e4f21dcc74d0e33ebfc08caa30e P  P         a   a   a   a             �"go.string.hdr.","                       go.string.","   �go.string.","   ,  �$go.string.hdr."!!"                       go.string."!!"   �go.string."!!"   !!  �"go.string.hdr."!"                       go.string."!"   �go.string."!"   !  �.go.string.hdr."android"                       &go.string."android"   �&go.string."android"   android  �Tgclocals·a95d0301643df1b330639fcf326ec36f 0  0           �          �Tgclocals·a4a72fe4111c0d730d77d6113711d8c8 0  0                   �(go.string.hdr."test"                        go.string."test"   � go.string."test"   
test  �Tgclocals·ac1513c540ef28dcd9fb2a42fdde591a                   �Tgclocals·c9451ec7b4e00af2b1e38fde82914877                  ��go.string.hdr."android darwin dragonfly freebsd linux nacl netbsd openbsd plan9 solaris windows "             Q          �go.string."android darwin dragonfly freebsd linux nacl netbsd openbsd plan9 solaris windows "   ��go.string."android darwin dragonfly freebsd linux nacl netbsd openbsd plan9 solaris windows " �  �android darwin dragonfly freebsd linux nacl netbsd openbsd plan9 solaris windows   �$"".hdr..gostring.1             �          ""..gostring.1   �""..gostring.1 �  �386 amd64 amd64p32 arm armbe arm64 arm64be ppc64 ppc64le mips mipsle mips64 mips64le mips64p32 mips64p32le ppc s390 s390x sparc sparc64   �Tgclocals·30fa7c694f0b53328be0204760229368               �    �Tgclocals·69c1753bd5f81501d95132d08af04464           �Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c      
        �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �dgo.string.hdr."architecture letter no longer used"             "          \go.string."architecture letter no longer used"   �\go.string."architecture letter no longer used" P  Farchitecture letter no longer used  �"go.string.hdr."?"                       go.string."?"   �go.string."?"   ?  �Tgclocals·11d28ee4a7546638afa514476454a63e (  (                 �Tgclocals·adb3347b296419e60da36d67f8b7ce43 (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Tgclocals·fce3d64185acee4a98aea2303545fc5c (  (                 �Tgclocals·f7309186bf9eeb0f8ece2eb16f2dc110 (  (                �^go.string.hdr."go/build: import reader looping"                       Vgo.string."go/build: import reader looping"   �Vgo.string."go/build: import reader looping" @  @go/build: import reader looping  �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Tgclocals·a1435607261436f22ba8c52b7acb6d2b (  (                 �Tgclocals·7e902992778eda5f91d29a3f0c115aee (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6             �Tgclocals·70b96bb4883c3816d291a08b355c816f @  @           �  �     0  0  �Tgclocals·28b6eb03a42390d78755fe1e234a72ea @  @                         �Tgclocals·8be1320446f57d096ee33ca6a889aca6 p  p   "           �      �             �      �      �Tgclocals·956d50cd930e9c0fc470cac7c8ba19b7 @  @   	                      �&go.string.hdr."lib"                       go.string."lib"   �go.string."lib"   lib  �$go.string.hdr.".a"                       go.string.".a"   �go.string.".a"   .a  �Tgclocals·d471303acc881ec3c678ddfbe4bb4911 `  `
                     R�� �� �� ��  ��  �Tgclocals·7be4bbacbfdb05fb3044e36c22b41e8b   
        �4go.string.hdr."/testdata/"             
          ,go.string."/testdata/"   �,go.string."/testdata/"    /testdata/  �2go.string.hdr."/testdata"             	          *go.string."/testdata"   �*go.string."/testdata"    /testdata  �2go.string.hdr."testdata/"             	          *go.string."testdata/"   �*go.string."testdata/"    testdata/  �0go.string.hdr."testdata"                       (go.string."testdata"   �(go.string."testdata"    testdata  �Tgclocals·63ba92e6c81d2d7bf2207e4076c8b23c      
        �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �(go.string.hdr."src/"                        go.string."src/"   � go.string."src/"   
src/  �,go.string.hdr."vendor"                       $go.string."vendor"   �$go.string."vendor"   vendor  �Tgclocals·68281ae9cb2c0df5f0c33d324dd29c1b �  �   (                 �     � �    ��     � 
    �       �T     �T      T     T       T      T   � 
     �Tgclocals·75ee4963a64d57666eac9d22b87e7339 �  �                                                 �Tgclocals·66499ec09befdf27c68e3e35878ba2c7 (  (                 �Tgclocals·7e902992778eda5f91d29a3f0c115aee (  (                �>""..gobytes.1   // �>""..gobytes.2   /* �>""..gobytes.3   */ �>""..gobytes.4   
 �>""..gobytes.5   // �>""..gobytes.6 �  � +-.,/0123456789=ABCDEFGHIJKLMNOPQRSTUVWXYZ_abcdefghijklmnopqrstuvwxyz:$@ �4go.string.hdr."darwin/386"             
          ,go.string."darwin/386"   �,go.string."darwin/386"    darwin/386  �8go.string.hdr."darwin/amd64"                       0go.string."darwin/amd64"   �0go.string."darwin/amd64"    darwin/amd64  �4go.string.hdr."darwin/arm"             
          ,go.string."darwin/arm"   �,go.string."darwin/arm"    darwin/arm  �8go.string.hdr."darwin/arm64"                       0go.string."darwin/arm64"   �0go.string."darwin/arm64"    darwin/arm64  �>go.string.hdr."dragonfly/amd64"                       6go.string."dragonfly/amd64"   �6go.string."dragonfly/amd64"     dragonfly/amd64  �6go.string.hdr."freebsd/386"                       .go.string."freebsd/386"   �.go.string."freebsd/386"    freebsd/386  �:go.string.hdr."freebsd/amd64"                       2go.string."freebsd/amd64"   �2go.string."freebsd/amd64"    freebsd/amd64  �6go.string.hdr."freebsd/arm"                       .go.string."freebsd/arm"   �.go.string."freebsd/arm"    freebsd/arm  �2go.string.hdr."linux/386"             	          *go.string."linux/386"   �*go.string."linux/386"    linux/386  �6go.string.hdr."linux/amd64"                       .go.string."linux/amd64"   �.go.string."linux/amd64"    linux/amd64  �2go.string.hdr."linux/arm"             	          *go.string."linux/arm"   �*go.string."linux/arm"    linux/arm  �6go.string.hdr."linux/arm64"                       .go.string."linux/arm64"   �.go.string."linux/arm64"    linux/arm64  �:go.string.hdr."linux/ppc64le"                       2go.string."linux/ppc64le"   �2go.string."linux/ppc64le"    linux/ppc64le  �6go.string.hdr."android/386"                       .go.string."android/386"   �.go.string."android/386"    android/386  �:go.string.hdr."android/amd64"                       2go.string."android/amd64"   �2go.string."android/amd64"    android/amd64  �6go.string.hdr."android/arm"                       .go.string."android/arm"   �.go.string."android/arm"    android/arm  �4go.string.hdr."netbsd/386"             
          ,go.string."netbsd/386"   �,go.string."netbsd/386"    netbsd/386  �8go.string.hdr."netbsd/amd64"                       0go.string."netbsd/amd64"   �0go.string."netbsd/amd64"    netbsd/amd64  �4go.string.hdr."netbsd/arm"             
          ,go.string."netbsd/arm"   �,go.string."netbsd/arm"    netbsd/arm  �6go.string.hdr."openbsd/386"                       .go.string."openbsd/386"   �.go.string."openbsd/386"    openbsd/386  �:go.string.hdr."openbsd/amd64"                       2go.string."openbsd/amd64"   �2go.string."openbsd/amd64"    openbsd/amd64  �:go.string.hdr."solaris/amd64"                       2go.string."solaris/amd64"   �2go.string."solaris/amd64"    solaris/amd64  �6go.string.hdr."windows/386"                       .go.string."windows/386"   �.go.string."windows/386"    windows/386  �:go.string.hdr."windows/amd64"                       2go.string."windows/amd64"   �2go.string."windows/amd64"    windows/amd64  �Hgo.string.hdr."pkg/tool/linux_amd64"                       @go.string."pkg/tool/linux_amd64"   �@go.string."pkg/tool/linux_amd64" 0  *pkg/tool/linux_amd64  �8go.string.hdr."syntax error"                       0go.string."syntax error"   �0go.string."syntax error"    syntax error  �Ngo.string.hdr."unexpected NUL in input"                       Fgo.string."unexpected NUL in input"   �Fgo.string."unexpected NUL in input" 0  0unexpected NUL in input  �Tgclocals·826f148c2b9ed682d2ed28d3c55a6368 (  (                 �Tgclocals·7d2d5fca80364273fb07d5820a76fef4           �<"".Default  �type."".Context   �<"".cgoEnabled  (type.map[string]bool   �:"".slashSlash  0type.[]uint8 0                         ""..gobytes.1   �:"".slashStar  0type.[]uint8 0                         ""..gobytes.2   �:"".starSlash  0type.[]uint8 0                         ""..gobytes.3   �:"".newline  0type.[]uint8 0                         ""..gobytes.4   �:"".slashslash  0type.[]uint8 0                         ""..gobytes.5   �:"".safeBytes  0type.[]uint8 0        I       I          ""..gobytes.6   �<"".knownOS  (type.map[string]bool   �<"".knownArch  (type.map[string]bool   �<"".ToolDir   type.string   �<"".errSyntax   type.error   �<"".errNUL   type.error   �""".statictmp_0062  @type.[2]string @                                  go.string."src"   �""".statictmp_0069  @type.[2]string @                                  go.string."src"   �""".statictmp_0086  �type.[6]string �                                                                                             "go.string."go1.1"      "go.string."go1.2"   @  "go.string."go1.3"   `  "go.string."go1.4"   �  "go.string."go1.5"   �  "go.string."go1.6"   �""".statictmp_0250  @type.[2]string @                                  go.string."src"   �""".statictmp_0257  @type.[2]string @                                  go.string."src"   �""".statictmp_0260  `type.[3]string @                                  go.string."src"   �""".statictmp_0267  `type.[3]string @                                  go.string."src"   �""".statictmp_0282  `type.[3]string @                                  go.string."src"   �""".statictmp_0291  `type.[3]string @                                  go.string."src"   �""".statictmp_0325  @type.[2]string @                                  go.string."src"   �""".statictmp_0328  @type.[2]string @                                  go.string."pkg"   �""".statictmp_0331  @type.[2]string @                                  go.string."bin"   �""".statictmp_0886  �type.[6]string �                                                                                                go.string."/"   `  go.string."lib"   �  go.string.".a"   �""".statictmp_0922  `type.[3]string `                                               @  $go.string."vendor"   �""".statictmp_0927  `type.[3]string @                                  $go.string."vendor"   �>"".initdone·  type.uint8   �""".statictmp_0939  �	Htype.[24]struct { a string; b bool } �        
                                            
                                                                                                                                    	                                            	                                                                                                                                    
                                            
                                                                                                                     0   ,go.string."darwin/386"   0  0go.string."darwin/amd64"   `  ,go.string."darwin/arm"   �  0go.string."darwin/arm64"   �  6go.string."dragonfly/amd64"   �  .go.string."freebsd/386"   �  2go.string."freebsd/amd64"   �  .go.string."freebsd/arm"   �  *go.string."linux/386"   �  .go.string."linux/amd64"   �  *go.string."linux/arm"   �  .go.string."linux/arm64"   �  2go.string."linux/ppc64le"   �  .go.string."android/386"   �  2go.string."android/amd64"   �  .go.string."android/arm"   �  ,go.string."netbsd/386"   �  0go.string."netbsd/amd64"   �  ,go.string."netbsd/arm"   �  .go.string."openbsd/386"   �  2go.string."openbsd/amd64"   �  2go.string."solaris/amd64"   �  .go.string."windows/386"   �  2go.string."windows/amd64"   �""".statictmp_0942  @type.[2]string @                                  @go.string."pkg/tool/linux_amd64"   �2"".(*Context).joinPath·f              ,"".(*Context).joinPath   �<"".(*Context).splitPathList·f              6"".(*Context).splitPathList   �4"".(*Context).isAbsPath·f              ."".(*Context).isAbsPath   �,"".(*Context).isDir·f              &"".(*Context).isDir   �4"".(*Context).hasSubdir·f              ."".(*Context).hasSubdir   �"".hasSubdir·f              "".hasSubdir   �0"".(*Context).readDir·f              *"".(*Context).readDir   �2"".(*Context).openFile·f              ,"".(*Context).openFile   �."".(*Context).isFile·f              ("".(*Context).isFile   �."".(*Context).gopath·f              ("".(*Context).gopath   �0"".(*Context).SrcDirs·f              *"".(*Context).SrcDirs   �("".defaultContext·f              """.defaultContext   �"".envOr·f              "".envOr   �4"".(*Package).IsCommand·f              ."".(*Package).IsCommand   �4"".(*Context).ImportDir·f              ."".(*Context).ImportDir   �0"".(*NoGoError).Error·f              *"".(*NoGoError).Error   �F"".(*MultiplePackageError).Error·f              @"".(*MultiplePackageError).Error   �"".nameExt·f              "".nameExt   �."".(*Context).Import·f              ("".(*Context).Import   � "".hasGoFiles·f              "".hasGoFiles   �."".findImportComment·f              ("".findImportComment   �0"".skipSpaceOrComment·f              *"".skipSpaceOrComment   �"".parseWord·f              "".parseWord   �4"".(*Context).MatchFile·f              ."".(*Context).MatchFile   �4"".(*Context).matchFile·f              ."".(*Context).matchFile   �$"".cleanImports·f              "".cleanImports   �"".Import·f              "".Import   �"".ImportDir·f              "".ImportDir   �8"".(*Context).shouldBuild·f              2"".(*Context).shouldBuild   �0"".(*Context).saveCgo·f              *"".(*Context).saveCgo   �$"".expandSrcDir·f              "".expandSrcDir   �""".safeCgoName·f              "".safeCgoName   �""".splitQuoted·f              "".splitQuoted   �,"".(*Context).match·f              &"".(*Context).match   �>"".(*Context).goodOSArchFile·f              8"".(*Context).goodOSArchFile   �"".init.1·f              "".init.1   �&"".IsLocalImport·f               "".IsLocalImport   �"".ArchChar·f              "".ArchChar   �"".isIdent·f              "".isIdent   �B"".(*importReader).syntaxError·f              <"".(*importReader).syntaxError   �<"".(*importReader).readByte·f              6"".(*importReader).readByte   �<"".(*importReader).peekByte·f              6"".(*importReader).peekByte   �<"".(*importReader).nextByte·f              6"".(*importReader).nextByte   �B"".(*importReader).readKeyword·f              <"".(*importReader).readKeyword   �>"".(*importReader).readIdent·f              8"".(*importReader).readIdent   �@"".(*importReader).readString·f              :"".(*importReader).readString   �@"".(*importReader).readImport·f              :"".(*importReader).readImport   �$"".readComments·f              "".readComments   �""".readImports·f              "".readImports   �:"".(*Context).Import.func1·f              4"".(*Context).Import.func1   �:"".(*Context).Import.func2·f              4"".(*Context).Import.func2   �:"".(*Context).Import.func3·f              4"".(*Context).Import.func3   �:"".(*Context).Import.func4·f              4"".(*Context).Import.func4   �"".init·f              "".init   �"runtime.gcbits.01    �0go.string.hdr."[]string"                       (go.string."[]string"   �(go.string."[]string"    []string  �type.[]string �  �              Ө�
                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  0go.string.hdr."[]string"   p  ,go.weak.type.*[]string   �  type.string   �:go.typelink.[]string	[]string              type.[]string   �Lgo.string.hdr."func(...string) string"                       Dgo.string."func(...string) string"   �Dgo.string."func(...string) string" 0  .func(...string) string  �6type.func(...string) string �  �              �l� 3                                                                                                           0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."func(...string) string"   p  Hgo.weak.type.*func(...string) string   �� 6type.func(...string) string   �� 6type.func(...string) string   �  type.[]string   �  type.string   �rgo.typelink.func(...string) string	func(...string) string              6type.func(...string) string   �Jgo.string.hdr."func(string) []string"                       Bgo.string."func(string) []string"   �Bgo.string."func(string) []string" 0  ,func(string) []string  �4type.func(string) []string �  �               �H� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Jgo.string.hdr."func(string) []string"   p  Fgo.weak.type.*func(string) []string   �� 4type.func(string) []string   �� 4type.func(string) []string   �  type.string   �  type.[]string   �ngo.typelink.func(string) []string	func(string) []string              4type.func(string) []string   �Bgo.string.hdr."func(string) bool"                       :go.string."func(string) bool"   �:go.string."func(string) bool" 0  $func(string) bool  �,type.func(string) bool �  �              *�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."func(string) bool"   p  >go.weak.type.*func(string) bool   �� ,type.func(string) bool   �� ,type.func(string) bool   �  type.string   �  type.bool   �^go.typelink.func(string) bool	func(string) bool              ,type.func(string) bool   �fgo.string.hdr."func(string, string) (string, bool)"             #          ^go.string."func(string, string) (string, bool)"   �^go.string."func(string, string) (string, bool)" P  Hfunc(string, string) (string, bool)  �Ptype.func(string, string) (string, bool) �  �              R�� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(string, string) (string, bool)"   p  bgo.weak.type.*func(string, string) (string, bool)   �� Ptype.func(string, string) (string, bool)   �� Ptype.func(string, string) (string, bool)   �  type.string   �  type.string   �  type.string   �  type.bool   ��go.typelink.func(string, string) (string, bool)	func(string, string) (string, bool)              Ptype.func(string, string) (string, bool)   �:go.string.hdr."[]os.FileInfo"                       2go.string."[]os.FileInfo"   �2go.string."[]os.FileInfo"    []os.FileInfo  �$type.[]os.FileInfo �  �              &�h                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."[]os.FileInfo"   p  6go.weak.type.*[]os.FileInfo   �   type.os.FileInfo   �Ngo.typelink.[]os.FileInfo	[]os.FileInfo              $type.[]os.FileInfo   �fgo.string.hdr."func(string) ([]os.FileInfo, error)"             #          ^go.string."func(string) ([]os.FileInfo, error)"   �^go.string."func(string) ([]os.FileInfo, error)" P  Hfunc(string) ([]os.FileInfo, error)  �Ptype.func(string) ([]os.FileInfo, error) �  �              ���� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(string) ([]os.FileInfo, error)"   p  bgo.weak.type.*func(string) ([]os.FileInfo, error)   �� Ptype.func(string) ([]os.FileInfo, error)   �� Ptype.func(string) ([]os.FileInfo, error)   �  type.string   �  $type.[]os.FileInfo   �  type.error   ��go.typelink.func(string) ([]os.FileInfo, error)	func(string) ([]os.FileInfo, error)              Ptype.func(string) ([]os.FileInfo, error)   �fgo.string.hdr."func(string) (io.ReadCloser, error)"             #          ^go.string."func(string) (io.ReadCloser, error)"   �^go.string."func(string) (io.ReadCloser, error)" P  Hfunc(string) (io.ReadCloser, error)  �Ptype.func(string) (io.ReadCloser, error) �  �              �?�p 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(string) (io.ReadCloser, error)"   p  bgo.weak.type.*func(string) (io.ReadCloser, error)   �� Ptype.func(string) (io.ReadCloser, error)   �� Ptype.func(string) (io.ReadCloser, error)   �  type.string   �  $type.io.ReadCloser   �  type.error   ��go.typelink.func(string) (io.ReadCloser, error)	func(string) (io.ReadCloser, error)              Ptype.func(string) (io.ReadCloser, error)   �.runtime.gcbits.554afa03   UJ� �:go.string.hdr."build.Context"                       2go.string."build.Context"   �2go.string."build.Context"    build.Context  �,go.string.hdr."GOROOT"                       $go.string."GOROOT"   �$go.string."GOROOT"   GOROOT  �4go.string.hdr."CgoEnabled"             
          ,go.string."CgoEnabled"   �,go.string."CgoEnabled"    CgoEnabled  �6go.string.hdr."UseAllFiles"                       .go.string."UseAllFiles"   �.go.string."UseAllFiles"    UseAllFiles  �0go.string.hdr."Compiler"                       (go.string."Compiler"   �(go.string."Compiler"    Compiler  �2go.string.hdr."BuildTags"             	          *go.string."BuildTags"   �*go.string."BuildTags"    BuildTags  �6go.string.hdr."ReleaseTags"                       .go.string."ReleaseTags"   �.go.string."ReleaseTags"    ReleaseTags  �:go.string.hdr."InstallSuffix"                       2go.string."InstallSuffix"   �2go.string."InstallSuffix"    InstallSuffix  �0go.string.hdr."JoinPath"                       (go.string."JoinPath"   �(go.string."JoinPath"    JoinPath  �:go.string.hdr."SplitPathList"                       2go.string."SplitPathList"   �2go.string."SplitPathList"    SplitPathList  �2go.string.hdr."IsAbsPath"             	          *go.string."IsAbsPath"   �*go.string."IsAbsPath"    IsAbsPath  �*go.string.hdr."IsDir"                       "go.string."IsDir"   �"go.string."IsDir"   IsDir  �2go.string.hdr."HasSubdir"             	          *go.string."HasSubdir"   �*go.string."HasSubdir"    HasSubdir  �.go.string.hdr."ReadDir"                       &go.string."ReadDir"   �&go.string."ReadDir"   ReadDir  �0go.string.hdr."OpenFile"                       (go.string."OpenFile"   �(go.string."OpenFile"    OpenFile  �.go.string.hdr."Context"                       &go.string."Context"   �&go.string."Context"   Context  �0go.string.hdr."go/build"                       (go.string."go/build"   �(go.string."go/build"    go/build  �"go.importpath."".                       (go.string."go/build"   �type."".Context  �  ��       �       ��G                                                                                                                                                                                                                      0                                       @                                       A                                       H                                       X                                       p                                       �                                       �                                       �                                       �                                       �                                       �                                       �                                       �                                               V0�  runtime.algarray   @  .runtime.gcbits.554afa03   P  :go.string.hdr."build.Context"   p   type.*"".Context   �� type."".Context   �  ,go.string.hdr."GOARCH"   �  type.string   �  (go.string.hdr."GOOS"   �  type.string   �  ,go.string.hdr."GOROOT"   �  type.string   �  ,go.string.hdr."GOPATH"   �  type.string   �  4go.string.hdr."CgoEnabled"   �  type.bool   �  6go.string.hdr."UseAllFiles"   �  type.bool   �  0go.string.hdr."Compiler"   �  type.string   �  2go.string.hdr."BuildTags"   �  type.[]string   �  6go.string.hdr."ReleaseTags"   �  type.[]string   �  :go.string.hdr."InstallSuffix"   �  type.string   �  0go.string.hdr."JoinPath"   �  6type.func(...string) string   �  :go.string.hdr."SplitPathList"   �  4type.func(string) []string   �  2go.string.hdr."IsAbsPath"   �	  ,type.func(string) bool   �	  *go.string.hdr."IsDir"   �	  ,type.func(string) bool   �
  2go.string.hdr."HasSubdir"   �
  Ptype.func(string, string) (string, bool)   �
  .go.string.hdr."ReadDir"   �  Ptype.func(string) ([]os.FileInfo, error)   �  0go.string.hdr."OpenFile"   �  Ptype.func(string) (io.ReadCloser, error)   `� type."".Context   �  .go.string.hdr."Context"   �  "go.importpath."".   �� type."".Context   �<go.string.hdr."*build.Context"                       4go.string."*build.Context"   �4go.string."*build.Context"    *build.Context  �Bgo.string.hdr."*build.ImportMode"                       :go.string."*build.ImportMode"   �:go.string."*build.ImportMode" 0  $*build.ImportMode  �&type.*"".ImportMode  �  �              U"l* 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."*build.ImportMode"   p  8go.weak.type.**"".ImportMode   �  $type."".ImportMode   �runtime.gcbits.      �@go.string.hdr."build.ImportMode"                       8go.string."build.ImportMode"   �8go.string."build.ImportMode" 0  "build.ImportMode  �4go.string.hdr."ImportMode"             
          ,go.string."ImportMode"   �,go.string."ImportMode"    ImportMode  �$type."".ImportMode  �  �               �~� �                                                                                0�  runtime.algarray   @  runtime.gcbits.   P  @go.string.hdr."build.ImportMode"   p  &type.*"".ImportMode   `� $type."".ImportMode   �  4go.string.hdr."ImportMode"   �  "go.importpath."".   �� $type."".ImportMode   �@go.string.hdr."[]token.Position"                       8go.string."[]token.Position"   �8go.string."[]token.Position" 0  "[]token.Position  �0type.[]go/token.Position �  �              f~��                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."[]token.Position"   p  Bgo.weak.type.*[]go/token.Position   �  ,type.go/token.Position   �`go.typelink.[]token.Position	[]go/token.Position              0type.[]go/token.Position   �.go.string.hdr."[]uint8"                       &go.string."[]uint8"   �&go.string."[]uint8"   []uint8  �type.[]uint8 �  �              �~.8                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  .go.string.hdr."[]uint8"   p  *go.weak.type.*[]uint8   �  type.uint8   �6go.typelink.[]uint8	[]uint8              type.[]uint8   �0go.string.hdr."[8]uint8"                       (go.string."[8]uint8"   �(go.string."[8]uint8"    [8]uint8  �type.[8]uint8 �  �               >�0� �                                                               0�  runtime.algarray   @  runtime.gcbits.   P  0go.string.hdr."[8]uint8"   p  ,go.weak.type.*[8]uint8   �  type.uint8   �  type.[]uint8   �:go.typelink.[8]uint8	[8]uint8              type.[8]uint8   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[8]string              (type..hash.[8]string   �,type..eqfunc.[8]string              $type..eq.[8]string   �&type..alg.[8]string                        0type..hashfunc.[8]string     ,type..eqfunc.[8]string   �&runtime.gcbits.5555   UU �2go.string.hdr."[8]string"             	          *go.string."[8]string"   �*go.string."[8]string"    [8]string  �type.[8]string �  ��       x       US�>                                                                0  &type..alg.[8]string   @  &runtime.gcbits.5555   P  2go.string.hdr."[8]string"   p  .go.weak.type.*[8]string   �  type.string   �  type.[]string   �>go.typelink.[8]string	[8]string              type.[8]string   �Dgo.string.hdr."[][]token.Position"                       <go.string."[][]token.Position"   �<go.string."[][]token.Position" 0  &[][]token.Position  �4type.[][]go/token.Position �  �              d� �                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."[][]token.Position"   p  Fgo.weak.type.*[][]go/token.Position   �  0type.[]go/token.Position   �hgo.typelink.[][]token.Position	[][]go/token.Position              4type.[][]go/token.Position   �*runtime.gcbits.499224   I�$ �Fgo.string.hdr."[8][]token.Position"                       >go.string."[8][]token.Position"   �>go.string."[8][]token.Position" 0  ([8][]token.Position  �6type.[8][]go/token.Position �  ��       �       ��s                                                                0�  runtime.algarray   @  *runtime.gcbits.499224   P  Fgo.string.hdr."[8][]token.Position"   p  Hgo.weak.type.*[8][]go/token.Position   �  0type.[]go/token.Position   �  4type.[][]go/token.Position   �lgo.typelink.[8][]token.Position	[8][]go/token.Position              6type.[8][]go/token.Position   �fgo.string.hdr."*map.bucket[string][]token.Position"             #          ^go.string."*map.bucket[string][]token.Position"   �^go.string."*map.bucket[string][]token.Position" P  H*map.bucket[string][]token.Position  �Vtype.*map.bucket[string][]go/token.Position �  �              ��9 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."*map.bucket[string][]token.Position"   p  hgo.weak.type.**map.bucket[string][]go/token.Position   �  Ttype.map.bucket[string][]go/token.Position   �6runtime.gcbits.aaaa92244902   ���$I �dgo.string.hdr."map.bucket[string][]token.Position"             "          \go.string."map.bucket[string][]token.Position"   �\go.string."map.bucket[string][]token.Position" P  Fmap.bucket[string][]token.Position  �.go.string.hdr."topbits"                       &go.string."topbits"   �&go.string."topbits"   topbits  �(go.string.hdr."keys"                        go.string."keys"   � go.string."keys"   
keys  �,go.string.hdr."values"                       $go.string."values"   �$go.string."values"   values  �0go.string.hdr."overflow"                       (go.string."overflow"   �(go.string."overflow"    overflow  �Ttype.map.bucket[string][]go/token.Position �  �P      P      RJ�x                                                                                                                                                                              �                                       H      0�  runtime.algarray   @  6runtime.gcbits.aaaa92244902   P  dgo.string.hdr."map.bucket[string][]token.Position"   p  fgo.weak.type.*map.bucket[string][]go/token.Position   �� Ttype.map.bucket[string][]go/token.Position   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  6type.[8][]go/token.Position   �  0go.string.hdr."overflow"   �  Vtype.*map.bucket[string][]go/token.Position   �"runtime.gcbits.2c   , �^go.string.hdr."map.hdr[string][]token.Position"                       Vgo.string."map.hdr[string][]token.Position"   �Vgo.string."map.hdr[string][]token.Position" @  @map.hdr[string][]token.Position  �*go.string.hdr."count"                       "go.string."count"   �"go.string."count"   count  �*go.string.hdr."flags"                       "go.string."flags"   �"go.string."flags"   flags  �"go.string.hdr."B"                       go.string."B"   �go.string."B"   B  �*go.string.hdr."hash0"                       "go.string."hash0"   �"go.string."hash0"   hash0  �.go.string.hdr."buckets"                       &go.string."buckets"   �&go.string."buckets"   buckets  �4go.string.hdr."oldbuckets"             
          ,go.string."oldbuckets"   �,go.string."oldbuckets"    oldbuckets  �2go.string.hdr."nevacuate"             	          *go.string."nevacuate"   �*go.string."nevacuate"    nevacuate  �Ntype.map.hdr[string][]go/token.Position �  �0       0       O��                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  ^go.string.hdr."map.hdr[string][]token.Position"   p  `go.weak.type.*map.hdr[string][]go/token.Position   �� Ntype.map.hdr[string][]go/token.Position   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  Vtype.*map.bucket[string][]go/token.Position   �  4go.string.hdr."oldbuckets"   �  Vtype.*map.bucket[string][]go/token.Position   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �Vgo.string.hdr."map[string][]token.Position"                       Ngo.string."map[string][]token.Position"   �Ngo.string."map[string][]token.Position" @  8map[string][]token.Position  �Ftype.map[string][]go/token.Position �  �              \�A	 5                                                                          P0�  runtime.algarray   @  "runtime.gcbits.01   P  Vgo.string.hdr."map[string][]token.Position"   p  Xgo.weak.type.*map[string][]go/token.Position   �  type.string   �  0type.[]go/token.Position   �  Ttype.map.bucket[string][]go/token.Position   �  Ntype.map.hdr[string][]go/token.Position   ��go.typelink.map[string][]token.Position	map[string][]go/token.Position              Ftype.map[string][]go/token.Position   �Rruntime.gcbits.5555a5942449922449924c2601   UU��$I�$I�L& �:go.string.hdr."build.Package"                       2go.string."build.Package"   �2go.string."build.Package"    build.Package  �&go.string.hdr."Dir"                       go.string."Dir"   �go.string."Dir"   Dir  �(go.string.hdr."Name"                        go.string."Name"   � go.string."Name"   
Name  �:go.string.hdr."ImportComment"                       2go.string."ImportComment"   �2go.string."ImportComment"    ImportComment  �&go.string.hdr."Doc"                       go.string."Doc"   �go.string."Doc"   Doc  �4go.string.hdr."ImportPath"             
          ,go.string."ImportPath"   �,go.string."ImportPath"    ImportPath  �(go.string.hdr."Root"                        go.string."Root"   � go.string."Root"   
Root  �.go.string.hdr."SrcRoot"                       &go.string."SrcRoot"   �&go.string."SrcRoot"   SrcRoot  �.go.string.hdr."PkgRoot"                       &go.string."PkgRoot"   �&go.string."PkgRoot"   PkgRoot  �:go.string.hdr."PkgTargetRoot"                       2go.string."PkgTargetRoot"   �2go.string."PkgTargetRoot"    PkgTargetRoot  �,go.string.hdr."BinDir"                       $go.string."BinDir"   �$go.string."BinDir"   BinDir  �,go.string.hdr."Goroot"                       $go.string."Goroot"   �$go.string."Goroot"   Goroot  �,go.string.hdr."PkgObj"                       $go.string."PkgObj"   �$go.string."PkgObj"   PkgObj  �.go.string.hdr."AllTags"                       &go.string."AllTags"   �&go.string."AllTags"   AllTags  �6go.string.hdr."ConflictDir"                       .go.string."ConflictDir"   �.go.string."ConflictDir"    ConflictDir  �.go.string.hdr."GoFiles"                       &go.string."GoFiles"   �&go.string."GoFiles"   GoFiles  �0go.string.hdr."CgoFiles"                       (go.string."CgoFiles"   �(go.string."CgoFiles"    CgoFiles  �<go.string.hdr."IgnoredGoFiles"                       4go.string."IgnoredGoFiles"   �4go.string."IgnoredGoFiles"    IgnoredGoFiles  �<go.string.hdr."InvalidGoFiles"                       4go.string."InvalidGoFiles"   �4go.string."InvalidGoFiles"    InvalidGoFiles  �,go.string.hdr."CFiles"                       $go.string."CFiles"   �$go.string."CFiles"   CFiles  �0go.string.hdr."CXXFiles"                       (go.string."CXXFiles"   �(go.string."CXXFiles"    CXXFiles  �,go.string.hdr."MFiles"                       $go.string."MFiles"   �$go.string."MFiles"   MFiles  �,go.string.hdr."HFiles"                       $go.string."HFiles"   �$go.string."HFiles"   HFiles  �,go.string.hdr."SFiles"                       $go.string."SFiles"   �$go.string."SFiles"   SFiles  �2go.string.hdr."SwigFiles"             	          *go.string."SwigFiles"   �*go.string."SwigFiles"    SwigFiles  �8go.string.hdr."SwigCXXFiles"                       0go.string."SwigCXXFiles"   �0go.string."SwigCXXFiles"    SwigCXXFiles  �2go.string.hdr."SysoFiles"             	          *go.string."SysoFiles"   �*go.string."SysoFiles"    SysoFiles  �2go.string.hdr."CgoCFLAGS"             	          *go.string."CgoCFLAGS"   �*go.string."CgoCFLAGS"    CgoCFLAGS  �6go.string.hdr."CgoCPPFLAGS"                       .go.string."CgoCPPFLAGS"   �.go.string."CgoCPPFLAGS"    CgoCPPFLAGS  �6go.string.hdr."CgoCXXFLAGS"                       .go.string."CgoCXXFLAGS"   �.go.string."CgoCXXFLAGS"    CgoCXXFLAGS  �4go.string.hdr."CgoLDFLAGS"             
          ,go.string."CgoLDFLAGS"   �,go.string."CgoLDFLAGS"    CgoLDFLAGS  �8go.string.hdr."CgoPkgConfig"                       0go.string."CgoPkgConfig"   �0go.string."CgoPkgConfig"    CgoPkgConfig  �.go.string.hdr."Imports"                       &go.string."Imports"   �&go.string."Imports"   Imports  �2go.string.hdr."ImportPos"             	          *go.string."ImportPos"   �*go.string."ImportPos"    ImportPos  �6go.string.hdr."TestGoFiles"                       .go.string."TestGoFiles"   �.go.string."TestGoFiles"    TestGoFiles  �6go.string.hdr."TestImports"                       .go.string."TestImports"   �.go.string."TestImports"    TestImports  �:go.string.hdr."TestImportPos"                       2go.string."TestImportPos"   �2go.string."TestImportPos"    TestImportPos  �8go.string.hdr."XTestGoFiles"                       0go.string."XTestGoFiles"   �0go.string."XTestGoFiles"    XTestGoFiles  �8go.string.hdr."XTestImports"                       0go.string."XTestImports"   �0go.string."XTestImports"    XTestImports  �<go.string.hdr."XTestImportPos"                       4go.string."XTestImportPos"   �4go.string."XTestImportPos"    XTestImportPos  �.go.string.hdr."Package"                       &go.string."Package"   �&go.string."Package"   Package  �type."".Package  �  �            �)Q�                                                 '       '                                                                                                                                                              0                                       @                                       P                                       `                                       p                                       �                                       �                                       �                                       �                                       �                                       �                                       �                                       �                                                                             (                                      @                                      X                                      p                                      �                                      �                                      �                                      �                                      �                                                                                                                   0                                      H                                      `                                      x                                      �                                      �                                      �                                      �                                      �                                      �                                                                                     �0�  runtime.algarray   @  Rruntime.gcbits.5555a5942449922449924c2601   P  :go.string.hdr."build.Package"   p   type.*"".Package   �� type."".Package   �  &go.string.hdr."Dir"   �  type.string   �  (go.string.hdr."Name"   �  type.string   �  :go.string.hdr."ImportComment"   �  type.string   �  &go.string.hdr."Doc"   �  type.string   �  4go.string.hdr."ImportPath"   �  type.string   �  (go.string.hdr."Root"   �  type.string   �  .go.string.hdr."SrcRoot"   �  type.string   �  .go.string.hdr."PkgRoot"   �  type.string   �  :go.string.hdr."PkgTargetRoot"   �  type.string   �  ,go.string.hdr."BinDir"   �  type.string   �  ,go.string.hdr."Goroot"   �  type.bool   �  ,go.string.hdr."PkgObj"   �  type.string   �  .go.string.hdr."AllTags"   �	  type.[]string   �	  6go.string.hdr."ConflictDir"   �	  type.string   �
  .go.string.hdr."GoFiles"   �
  type.[]string   �
  0go.string.hdr."CgoFiles"   �  type.[]string   �  <go.string.hdr."IgnoredGoFiles"   �  type.[]string   �  <go.string.hdr."InvalidGoFiles"   �  type.[]string   �  ,go.string.hdr."CFiles"   �  type.[]string   �  0go.string.hdr."CXXFiles"   �  type.[]string   �  ,go.string.hdr."MFiles"   �  type.[]string   �  ,go.string.hdr."HFiles"   �  type.[]string   �  ,go.string.hdr."SFiles"   �  type.[]string   �  2go.string.hdr."SwigFiles"   �  type.[]string   �  8go.string.hdr."SwigCXXFiles"   �  type.[]string   �  2go.string.hdr."SysoFiles"   �  type.[]string   �  2go.string.hdr."CgoCFLAGS"   �  type.[]string   �  6go.string.hdr."CgoCPPFLAGS"   �  type.[]string   �  6go.string.hdr."CgoCXXFLAGS"   �  type.[]string   �  4go.string.hdr."CgoLDFLAGS"   �  type.[]string   �  8go.string.hdr."CgoPkgConfig"   �  type.[]string   �  .go.string.hdr."Imports"   �  type.[]string   �  2go.string.hdr."ImportPos"   �  Ftype.map[string][]go/token.Position   �  6go.string.hdr."TestGoFiles"   �  type.[]string   �  6go.string.hdr."TestImports"   �  type.[]string   �  :go.string.hdr."TestImportPos"   �  Ftype.map[string][]go/token.Position   �  8go.string.hdr."XTestGoFiles"   �  type.[]string   �  8go.string.hdr."XTestImports"   �  type.[]string   �  <go.string.hdr."XTestImportPos"   �  Ftype.map[string][]go/token.Position   `� type."".Package   �  .go.string.hdr."Package"   �  "go.importpath."".   �� type."".Package   �<go.string.hdr."*build.Package"                       4go.string."*build.Package"   �4go.string."*build.Package"    *build.Package  �Rgo.string.hdr."func(*build.Package) bool"                       Jgo.string."func(*build.Package) bool"   �Jgo.string."func(*build.Package) bool" @  4func(*build.Package) bool  �6type.func(*"".Package) bool �  �              �s�t 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func(*build.Package) bool"   p  Hgo.weak.type.*func(*"".Package) bool   �� 6type.func(*"".Package) bool   �� 6type.func(*"".Package) bool   �   type.*"".Package   �  type.bool   �xgo.typelink.func(*build.Package) bool	func(*"".Package) bool              6type.func(*"".Package) bool   �2go.string.hdr."IsCommand"             	          *go.string."IsCommand"   �*go.string."IsCommand"    IsCommand  �6go.string.hdr."func() bool"                       .go.string."func() bool"   �.go.string."func() bool"    func() bool  � type.func() bool �  �              T�x 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."func() bool"   p  2go.weak.type.*func() bool   ��  type.func() bool   ��  type.func() bool   �  type.bool   �Fgo.typelink.func() bool	func() bool               type.func() bool   � type.*"".Package  �  �              �)�� 6                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."*build.Package"   p  2go.weak.type.**"".Package   �  type."".Package   `�  type.*"".Package   ��  type.*"".Package   �  2go.string.hdr."IsCommand"   �   type.func() bool   �  6type.func(*"".Package) bool   �  ."".(*Package).IsCommand   �  ."".(*Package).IsCommand   ��go.string.hdr."func(*build.Context, string, string, build.ImportMode) (*build.Package, error)"             N          �go.string."func(*build.Context, string, string, build.ImportMode) (*build.Package, error)"   ��go.string."func(*build.Context, string, string, build.ImportMode) (*build.Package, error)" �  �func(*build.Context, string, string, build.ImportMode) (*build.Package, error)  ��type.func(*"".Context, string, string, "".ImportMode) (*"".Package, error) �  �              L� 3                                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, string, build.ImportMode) (*build.Package, error)"   p  �go.weak.type.*func(*"".Context, string, string, "".ImportMode) (*"".Package, error)   �� �type.func(*"".Context, string, string, "".ImportMode) (*"".Package, error)   �� �type.func(*"".Context, string, string, "".ImportMode) (*"".Package, error)   �   type.*"".Context   �  type.string   �  type.string   �  $type."".ImportMode   �   type.*"".Package   �  type.error   ��go.typelink.func(*build.Context, string, string, build.ImportMode) (*build.Package, error)	func(*"".Context, string, string, "".ImportMode) (*"".Package, error)              �type.func(*"".Context, string, string, "".ImportMode) (*"".Package, error)   ��go.string.hdr."func(*build.Context, string, build.ImportMode) (*build.Package, error)"             F          �go.string."func(*build.Context, string, build.ImportMode) (*build.Package, error)"   ��go.string."func(*build.Context, string, build.ImportMode) (*build.Package, error)" �  �func(*build.Context, string, build.ImportMode) (*build.Package, error)  ��type.func(*"".Context, string, "".ImportMode) (*"".Package, error) �  �              �; 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, build.ImportMode) (*build.Package, error)"   p  �go.weak.type.*func(*"".Context, string, "".ImportMode) (*"".Package, error)   �� �type.func(*"".Context, string, "".ImportMode) (*"".Package, error)   �� �type.func(*"".Context, string, "".ImportMode) (*"".Package, error)   �   type.*"".Context   �  type.string   �  $type."".ImportMode   �   type.*"".Package   �  type.error   ��go.typelink.func(*build.Context, string, build.ImportMode) (*build.Package, error)	func(*"".Context, string, "".ImportMode) (*"".Package, error)              �type.func(*"".Context, string, "".ImportMode) (*"".Package, error)   ��go.string.hdr."func(*build.Context, string, string) (bool, error)"             2          |go.string."func(*build.Context, string, string) (bool, error)"   �|go.string."func(*build.Context, string, string) (bool, error)" p  ffunc(*build.Context, string, string) (bool, error)  �htype.func(*"".Context, string, string) (bool, error) �  �              ��c 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, string) (bool, error)"   p  zgo.weak.type.*func(*"".Context, string, string) (bool, error)   �� htype.func(*"".Context, string, string) (bool, error)   �� htype.func(*"".Context, string, string) (bool, error)   �   type.*"".Context   �  type.string   �  type.string   �  type.bool   �  type.error   ��go.typelink.func(*build.Context, string, string) (bool, error)	func(*"".Context, string, string) (bool, error)              htype.func(*"".Context, string, string) (bool, error)   �Zgo.string.hdr."func(*build.Context) []string"                       Rgo.string."func(*build.Context) []string"   �Rgo.string."func(*build.Context) []string" @  <func(*build.Context) []string  �>type.func(*"".Context) []string �  �              � 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."func(*build.Context) []string"   p  Pgo.weak.type.*func(*"".Context) []string   �� >type.func(*"".Context) []string   �� >type.func(*"".Context) []string   �   type.*"".Context   �  type.[]string   ��go.typelink.func(*build.Context) []string	func(*"".Context) []string              >type.func(*"".Context) []string   �,go.string.hdr."[]bool"                       $go.string."[]bool"   �$go.string."[]bool"   []bool  �type.[]bool �  �              ���                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  ,go.string.hdr."[]bool"   p  (go.weak.type.*[]bool   �  type.bool   �2go.typelink.[]bool	[]bool              type.[]bool   �.go.string.hdr."[8]bool"                       &go.string."[8]bool"   �&go.string."[8]bool"   [8]bool  �type.[8]bool �  �               s�5 �                                                               0�  runtime.algarray   @  runtime.gcbits.   P  .go.string.hdr."[8]bool"   p  *go.weak.type.*[8]bool   �  type.bool   �  type.[]bool   �6go.typelink.[8]bool	[8]bool              type.[8]bool   �Ngo.string.hdr."*map.bucket[string]bool"                       Fgo.string."*map.bucket[string]bool"   �Fgo.string."*map.bucket[string]bool" 0  0*map.bucket[string]bool  �8type.*map.bucket[string]bool �  �              �[�E 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."*map.bucket[string]bool"   p  Jgo.weak.type.**map.bucket[string]bool   �  6type.map.bucket[string]bool   �*runtime.gcbits.aaaa04   �� �Lgo.string.hdr."map.bucket[string]bool"                       Dgo.string."map.bucket[string]bool"   �Dgo.string."map.bucket[string]bool" 0  .map.bucket[string]bool  �6type.map.bucket[string]bool �  ��       �       2aB�                                                                                                                                                                              �                                       �       0�  runtime.algarray   @  *runtime.gcbits.aaaa04   P  Lgo.string.hdr."map.bucket[string]bool"   p  Hgo.weak.type.*map.bucket[string]bool   �� 6type.map.bucket[string]bool   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  type.[8]bool   �  0go.string.hdr."overflow"   �  8type.*map.bucket[string]bool   �Fgo.string.hdr."map.hdr[string]bool"                       >go.string."map.hdr[string]bool"   �>go.string."map.hdr[string]bool" 0  (map.hdr[string]bool  �0type.map.hdr[string]bool �  �0       0       3�(                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Fgo.string.hdr."map.hdr[string]bool"   p  Bgo.weak.type.*map.hdr[string]bool   �� 0type.map.hdr[string]bool   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  8type.*map.bucket[string]bool   �  4go.string.hdr."oldbuckets"   �  8type.*map.bucket[string]bool   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �>go.string.hdr."map[string]bool"                       6go.string."map[string]bool"   �6go.string."map[string]bool"     map[string]bool  �(type.map[string]bool �  �              �� 5                                                                          � 0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."map[string]bool"   p  :go.weak.type.*map[string]bool   �  type.string   �  type.bool   �  6type.map.bucket[string]bool   �  0type.map.hdr[string]bool   �Vgo.typelink.map[string]bool	map[string]bool              (type.map[string]bool   ��go.string.hdr."func(*build.Context, string, map[string]bool) bool"             2          |go.string."func(*build.Context, string, map[string]bool) bool"   �|go.string."func(*build.Context, string, map[string]bool) bool" p  ffunc(*build.Context, string, map[string]bool) bool  �htype.func(*"".Context, string, map[string]bool) bool �  �              �! 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, map[string]bool) bool"   p  zgo.weak.type.*func(*"".Context, string, map[string]bool) bool   �� htype.func(*"".Context, string, map[string]bool) bool   �� htype.func(*"".Context, string, map[string]bool) bool   �   type.*"".Context   �  type.string   �  (type.map[string]bool   �  type.bool   ��go.typelink.func(*build.Context, string, map[string]bool) bool	func(*"".Context, string, map[string]bool) bool              htype.func(*"".Context, string, map[string]bool) bool   ��go.string.hdr."func(*build.Context, string, string) (string, bool)"             3          ~go.string."func(*build.Context, string, string) (string, bool)"   �~go.string."func(*build.Context, string, string) (string, bool)" p  hfunc(*build.Context, string, string) (string, bool)  �jtype.func(*"".Context, string, string) (string, bool) �  �              -"=� 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, string) (string, bool)"   p  |go.weak.type.*func(*"".Context, string, string) (string, bool)   �� jtype.func(*"".Context, string, string) (string, bool)   �� jtype.func(*"".Context, string, string) (string, bool)   �   type.*"".Context   �  type.string   �  type.string   �  type.string   �  type.bool   ��go.typelink.func(*build.Context, string, string) (string, bool)	func(*"".Context, string, string) (string, bool)              jtype.func(*"".Context, string, string) (string, bool)   �bgo.string.hdr."func(*build.Context, string) bool"             !          Zgo.string."func(*build.Context, string) bool"   �Zgo.string."func(*build.Context, string) bool" P  Dfunc(*build.Context, string) bool  �Ftype.func(*"".Context, string) bool �  �              �`�� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*build.Context, string) bool"   p  Xgo.weak.type.*func(*"".Context, string) bool   �� Ftype.func(*"".Context, string) bool   �� Ftype.func(*"".Context, string) bool   �   type.*"".Context   �  type.string   �  type.bool   ��go.typelink.func(*build.Context, string) bool	func(*"".Context, string) bool              Ftype.func(*"".Context, string) bool   �lgo.string.hdr."func(*build.Context, ...string) string"             &          dgo.string."func(*build.Context, ...string) string"   �dgo.string."func(*build.Context, ...string) string" P  Nfunc(*build.Context, ...string) string  �Ptype.func(*"".Context, ...string) string �  �              �I�+ 3                                                                                                                   0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(*build.Context, ...string) string"   p  bgo.weak.type.*func(*"".Context, ...string) string   �� Ptype.func(*"".Context, ...string) string   �� Ptype.func(*"".Context, ...string) string   �   type.*"".Context   �  type.[]string   �  type.string   ��go.typelink.func(*build.Context, ...string) string	func(*"".Context, ...string) string              Ptype.func(*"".Context, ...string) string   ��go.string.hdr."func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)"             Z          �go.string."func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)"   ��go.string."func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)" �  �func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)  ��type.func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error) �  �              �� 3                                                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)"   p  �go.weak.type.*func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)   �� �type.func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)   �� �type.func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)   �   type.*"".Context   �  type.string   �  type.string   �  type.bool   �  (type.map[string]bool   �  type.bool   �  type.[]uint8   �  type.string   �  type.error   ��go.typelink.func(*build.Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)	func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)              �type.func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)   ��go.string.hdr."func(*build.Context, string) (io.ReadCloser, error)"             3          ~go.string."func(*build.Context, string) (io.ReadCloser, error)"   �~go.string."func(*build.Context, string) (io.ReadCloser, error)" p  hfunc(*build.Context, string) (io.ReadCloser, error)  �jtype.func(*"".Context, string) (io.ReadCloser, error) �  �              �>�� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string) (io.ReadCloser, error)"   p  |go.weak.type.*func(*"".Context, string) (io.ReadCloser, error)   �� jtype.func(*"".Context, string) (io.ReadCloser, error)   �� jtype.func(*"".Context, string) (io.ReadCloser, error)   �   type.*"".Context   �  type.string   �  $type.io.ReadCloser   �  type.error   ��go.typelink.func(*build.Context, string) (io.ReadCloser, error)	func(*"".Context, string) (io.ReadCloser, error)              jtype.func(*"".Context, string) (io.ReadCloser, error)   ��go.string.hdr."func(*build.Context, string) ([]os.FileInfo, error)"             3          ~go.string."func(*build.Context, string) ([]os.FileInfo, error)"   �~go.string."func(*build.Context, string) ([]os.FileInfo, error)" p  hfunc(*build.Context, string) ([]os.FileInfo, error)  �jtype.func(*"".Context, string) ([]os.FileInfo, error) �  �              �nJ 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string) ([]os.FileInfo, error)"   p  |go.weak.type.*func(*"".Context, string) ([]os.FileInfo, error)   �� jtype.func(*"".Context, string) ([]os.FileInfo, error)   �� jtype.func(*"".Context, string) ([]os.FileInfo, error)   �   type.*"".Context   �  type.string   �  $type.[]os.FileInfo   �  type.error   ��go.typelink.func(*build.Context, string) ([]os.FileInfo, error)	func(*"".Context, string) ([]os.FileInfo, error)              jtype.func(*"".Context, string) ([]os.FileInfo, error)   ��go.string.hdr."func(*build.Context, string, *build.Package, *ast.CommentGroup) error"             E          �go.string."func(*build.Context, string, *build.Package, *ast.CommentGroup) error"   ��go.string."func(*build.Context, string, *build.Package, *ast.CommentGroup) error" �  �func(*build.Context, string, *build.Package, *ast.CommentGroup) error  ��type.func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error �  �               ��� 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, string, *build.Package, *ast.CommentGroup) error"   p  �go.weak.type.*func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error   �� �type.func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error   �� �type.func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error   �   type.*"".Context   �  type.string   �   type.*"".Package   �  2type.*go/ast.CommentGroup   �  type.error   ��go.typelink.func(*build.Context, string, *build.Package, *ast.CommentGroup) error	func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error              �type.func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error   ��go.string.hdr."func(*build.Context, []uint8, map[string]bool) bool"             3          ~go.string."func(*build.Context, []uint8, map[string]bool) bool"   �~go.string."func(*build.Context, []uint8, map[string]bool) bool" p  hfunc(*build.Context, []uint8, map[string]bool) bool  �jtype.func(*"".Context, []uint8, map[string]bool) bool �  �              cMo� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*build.Context, []uint8, map[string]bool) bool"   p  |go.weak.type.*func(*"".Context, []uint8, map[string]bool) bool   �� jtype.func(*"".Context, []uint8, map[string]bool) bool   �� jtype.func(*"".Context, []uint8, map[string]bool) bool   �   type.*"".Context   �  type.[]uint8   �  (type.map[string]bool   �  type.bool   ��go.typelink.func(*build.Context, []uint8, map[string]bool) bool	func(*"".Context, []uint8, map[string]bool) bool              jtype.func(*"".Context, []uint8, map[string]bool) bool   �jgo.string.hdr."func(*build.Context, string) []string"             %          bgo.string."func(*build.Context, string) []string"   �bgo.string."func(*build.Context, string) []string" P  Lfunc(*build.Context, string) []string  �Ntype.func(*"".Context, string) []string �  �              ,��u 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(*build.Context, string) []string"   p  `go.weak.type.*func(*"".Context, string) []string   �� Ntype.func(*"".Context, string) []string   �� Ntype.func(*"".Context, string) []string   �   type.*"".Context   �  type.string   �  type.[]string   ��go.typelink.func(*build.Context, string) []string	func(*"".Context, string) []string              Ntype.func(*"".Context, string) []string   �,go.string.hdr."Import"                       $go.string."Import"   �$go.string."Import"   Import  ��go.string.hdr."func(string, string, build.ImportMode) (*build.Package, error)"             >          �go.string."func(string, string, build.ImportMode) (*build.Package, error)"   ��go.string."func(string, string, build.ImportMode) (*build.Package, error)" �  ~func(string, string, build.ImportMode) (*build.Package, error)  �ztype.func(string, string, "".ImportMode) (*"".Package, error) �  �              ���> 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(string, string, build.ImportMode) (*build.Package, error)"   p  �go.weak.type.*func(string, string, "".ImportMode) (*"".Package, error)   �� ztype.func(string, string, "".ImportMode) (*"".Package, error)   �� ztype.func(string, string, "".ImportMode) (*"".Package, error)   �  type.string   �  type.string   �  $type."".ImportMode   �   type.*"".Package   �  type.error   ��go.typelink.func(string, string, build.ImportMode) (*build.Package, error)	func(string, string, "".ImportMode) (*"".Package, error)              ztype.func(string, string, "".ImportMode) (*"".Package, error)   �2go.string.hdr."ImportDir"             	          *go.string."ImportDir"   �*go.string."ImportDir"    ImportDir  ��go.string.hdr."func(string, build.ImportMode) (*build.Package, error)"             6          �go.string."func(string, build.ImportMode) (*build.Package, error)"   ��go.string."func(string, build.ImportMode) (*build.Package, error)" p  nfunc(string, build.ImportMode) (*build.Package, error)  �jtype.func(string, "".ImportMode) (*"".Package, error) �  �              �;5j 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(string, build.ImportMode) (*build.Package, error)"   p  |go.weak.type.*func(string, "".ImportMode) (*"".Package, error)   �� jtype.func(string, "".ImportMode) (*"".Package, error)   �� jtype.func(string, "".ImportMode) (*"".Package, error)   �  type.string   �  $type."".ImportMode   �   type.*"".Package   �  type.error   ��go.typelink.func(string, build.ImportMode) (*build.Package, error)	func(string, "".ImportMode) (*"".Package, error)              jtype.func(string, "".ImportMode) (*"".Package, error)   �2go.string.hdr."MatchFile"             	          *go.string."MatchFile"   �*go.string."MatchFile"    MatchFile  �dgo.string.hdr."func(string, string) (bool, error)"             "          \go.string."func(string, string) (bool, error)"   �\go.string."func(string, string) (bool, error)" P  Ffunc(string, string) (bool, error)  �Ntype.func(string, string) (bool, error) �  �              B�7# 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  dgo.string.hdr."func(string, string) (bool, error)"   p  `go.weak.type.*func(string, string) (bool, error)   �� Ntype.func(string, string) (bool, error)   �� Ntype.func(string, string) (bool, error)   �  type.string   �  type.string   �  type.bool   �  type.error   ��go.typelink.func(string, string) (bool, error)	func(string, string) (bool, error)              Ntype.func(string, string) (bool, error)   �.go.string.hdr."SrcDirs"                       &go.string."SrcDirs"   �&go.string."SrcDirs"   SrcDirs  �>go.string.hdr."func() []string"                       6go.string."func() []string"   �6go.string."func() []string"     func() []string  �(type.func() []string �  �              ���� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."func() []string"   p  :go.weak.type.*func() []string   �� (type.func() []string   �� (type.func() []string   �  type.[]string   �Vgo.typelink.func() []string	func() []string              (type.func() []string   �<go.string.hdr."goodOSArchFile"                       4go.string."goodOSArchFile"   �4go.string."goodOSArchFile"    goodOSArchFile  �dgo.string.hdr."func(string, map[string]bool) bool"             "          \go.string."func(string, map[string]bool) bool"   �\go.string."func(string, map[string]bool) bool" P  Ffunc(string, map[string]bool) bool  �Ntype.func(string, map[string]bool) bool �  �              I��  3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  dgo.string.hdr."func(string, map[string]bool) bool"   p  `go.weak.type.*func(string, map[string]bool) bool   �� Ntype.func(string, map[string]bool) bool   �� Ntype.func(string, map[string]bool) bool   �  type.string   �  (type.map[string]bool   �  type.bool   ��go.typelink.func(string, map[string]bool) bool	func(string, map[string]bool) bool              Ntype.func(string, map[string]bool) bool   �,go.string.hdr."gopath"                       $go.string."gopath"   �$go.string."gopath"   gopath  �2go.string.hdr."hasSubdir"             	          *go.string."hasSubdir"   �*go.string."hasSubdir"    hasSubdir  �2go.string.hdr."isAbsPath"             	          *go.string."isAbsPath"   �*go.string."isAbsPath"    isAbsPath  �*go.string.hdr."isDir"                       "go.string."isDir"   �"go.string."isDir"   isDir  �,go.string.hdr."isFile"                       $go.string."isFile"   �$go.string."isFile"   isFile  �0go.string.hdr."joinPath"                       (go.string."joinPath"   �(go.string."joinPath"    joinPath  �*go.string.hdr."match"                       "go.string."match"   �"go.string."match"   match  �2go.string.hdr."matchFile"             	          *go.string."matchFile"   �*go.string."matchFile"    matchFile  ��go.string.hdr."func(string, string, bool, map[string]bool) (bool, []uint8, string, error)"             J          �go.string."func(string, string, bool, map[string]bool) (bool, []uint8, string, error)"   ��go.string."func(string, string, bool, map[string]bool) (bool, []uint8, string, error)" �  �func(string, string, bool, map[string]bool) (bool, []uint8, string, error)  ��type.func(string, string, bool, map[string]bool) (bool, []uint8, string, error) �  �              ئ� 3                                                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(string, string, bool, map[string]bool) (bool, []uint8, string, error)"   p  �go.weak.type.*func(string, string, bool, map[string]bool) (bool, []uint8, string, error)   �� �type.func(string, string, bool, map[string]bool) (bool, []uint8, string, error)   �� �type.func(string, string, bool, map[string]bool) (bool, []uint8, string, error)   �  type.string   �  type.string   �  type.bool   �  (type.map[string]bool   �  type.bool   �  type.[]uint8   �  type.string   �  type.error   ��go.typelink.func(string, string, bool, map[string]bool) (bool, []uint8, string, error)	func(string, string, bool, map[string]bool) (bool, []uint8, string, error)              �type.func(string, string, bool, map[string]bool) (bool, []uint8, string, error)   �0go.string.hdr."openFile"                       (go.string."openFile"   �(go.string."openFile"    openFile  �.go.string.hdr."readDir"                       &go.string."readDir"   �&go.string."readDir"   readDir  �.go.string.hdr."saveCgo"                       &go.string."saveCgo"   �&go.string."saveCgo"   saveCgo  ��go.string.hdr."func(string, *build.Package, *ast.CommentGroup) error"             5          �go.string."func(string, *build.Package, *ast.CommentGroup) error"   ��go.string."func(string, *build.Package, *ast.CommentGroup) error" p  lfunc(string, *build.Package, *ast.CommentGroup) error  �ttype.func(string, *"".Package, *go/ast.CommentGroup) error �  �              ��T 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(string, *build.Package, *ast.CommentGroup) error"   p  �go.weak.type.*func(string, *"".Package, *go/ast.CommentGroup) error   �� ttype.func(string, *"".Package, *go/ast.CommentGroup) error   �� ttype.func(string, *"".Package, *go/ast.CommentGroup) error   �  type.string   �   type.*"".Package   �  2type.*go/ast.CommentGroup   �  type.error   ��go.typelink.func(string, *build.Package, *ast.CommentGroup) error	func(string, *"".Package, *go/ast.CommentGroup) error              ttype.func(string, *"".Package, *go/ast.CommentGroup) error   �6go.string.hdr."shouldBuild"                       .go.string."shouldBuild"   �.go.string."shouldBuild"    shouldBuild  �fgo.string.hdr."func([]uint8, map[string]bool) bool"             #          ^go.string."func([]uint8, map[string]bool) bool"   �^go.string."func([]uint8, map[string]bool) bool" P  Hfunc([]uint8, map[string]bool) bool  �Ptype.func([]uint8, map[string]bool) bool �  �              �!�; 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func([]uint8, map[string]bool) bool"   p  bgo.weak.type.*func([]uint8, map[string]bool) bool   �� Ptype.func([]uint8, map[string]bool) bool   �� Ptype.func([]uint8, map[string]bool) bool   �  type.[]uint8   �  (type.map[string]bool   �  type.bool   ��go.typelink.func([]uint8, map[string]bool) bool	func([]uint8, map[string]bool) bool              Ptype.func([]uint8, map[string]bool) bool   �:go.string.hdr."splitPathList"                       2go.string."splitPathList"   �2go.string."splitPathList"    splitPathList  � type.*"".Context  �  �              �V�I 6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."*build.Context"   p  2go.weak.type.**"".Context   �  type."".Context   `�  type.*"".Context   ��  type.*"".Context   �  ,go.string.hdr."Import"   �  ztype.func(string, string, "".ImportMode) (*"".Package, error)   �  �type.func(*"".Context, string, string, "".ImportMode) (*"".Package, error)   �  ("".(*Context).Import   �  ("".(*Context).Import   �  2go.string.hdr."ImportDir"   �  jtype.func(string, "".ImportMode) (*"".Package, error)   �  �type.func(*"".Context, string, "".ImportMode) (*"".Package, error)   �  ."".(*Context).ImportDir   �  ."".(*Context).ImportDir   �  2go.string.hdr."MatchFile"   �  Ntype.func(string, string) (bool, error)   �  htype.func(*"".Context, string, string) (bool, error)   �  ."".(*Context).MatchFile   �  ."".(*Context).MatchFile   �  .go.string.hdr."SrcDirs"   �  (type.func() []string   �  >type.func(*"".Context) []string   �  *"".(*Context).SrcDirs   �  *"".(*Context).SrcDirs   �  <go.string.hdr."goodOSArchFile"   �  "go.importpath."".   �  Ntype.func(string, map[string]bool) bool   �  htype.func(*"".Context, string, map[string]bool) bool   �  8"".(*Context).goodOSArchFile   �  8"".(*Context).goodOSArchFile   �  ,go.string.hdr."gopath"   �  "go.importpath."".   �  (type.func() []string   �  >type.func(*"".Context) []string   �  ("".(*Context).gopath   �  ("".(*Context).gopath   �  2go.string.hdr."hasSubdir"   �  "go.importpath."".   �  Ptype.func(string, string) (string, bool)   �  jtype.func(*"".Context, string, string) (string, bool)   �  ."".(*Context).hasSubdir   �  ."".(*Context).hasSubdir   �  2go.string.hdr."isAbsPath"   �  "go.importpath."".   �  ,type.func(string) bool   �  Ftype.func(*"".Context, string) bool   �  ."".(*Context).isAbsPath   �  ."".(*Context).isAbsPath   �  *go.string.hdr."isDir"   �  "go.importpath."".   �  ,type.func(string) bool   �  Ftype.func(*"".Context, string) bool   �  &"".(*Context).isDir   �  &"".(*Context).isDir   �  ,go.string.hdr."isFile"   �  "go.importpath."".   �  ,type.func(string) bool   �  Ftype.func(*"".Context, string) bool   �	  ("".(*Context).isFile   �	  ("".(*Context).isFile   �	  0go.string.hdr."joinPath"   �	  "go.importpath."".   �	  6type.func(...string) string   �	  Ptype.func(*"".Context, ...string) string   �	  ,"".(*Context).joinPath   �	  ,"".(*Context).joinPath   �
  *go.string.hdr."match"   �
  "go.importpath."".   �
  Ntype.func(string, map[string]bool) bool   �
  htype.func(*"".Context, string, map[string]bool) bool   �
  &"".(*Context).match   �
  &"".(*Context).match   �
  2go.string.hdr."matchFile"   �
  "go.importpath."".   �  �type.func(string, string, bool, map[string]bool) (bool, []uint8, string, error)   �  �type.func(*"".Context, string, string, bool, map[string]bool) (bool, []uint8, string, error)   �  ."".(*Context).matchFile   �  ."".(*Context).matchFile   �  0go.string.hdr."openFile"   �  "go.importpath."".   �  Ptype.func(string) (io.ReadCloser, error)   �  jtype.func(*"".Context, string) (io.ReadCloser, error)   �  ,"".(*Context).openFile   �  ,"".(*Context).openFile   �  .go.string.hdr."readDir"   �  "go.importpath."".   �  Ptype.func(string) ([]os.FileInfo, error)   �  jtype.func(*"".Context, string) ([]os.FileInfo, error)   �  *"".(*Context).readDir   �  *"".(*Context).readDir   �  .go.string.hdr."saveCgo"   �  "go.importpath."".   �  ttype.func(string, *"".Package, *go/ast.CommentGroup) error   �  �type.func(*"".Context, string, *"".Package, *go/ast.CommentGroup) error   �  *"".(*Context).saveCgo   �  *"".(*Context).saveCgo   �  6go.string.hdr."shouldBuild"   �  "go.importpath."".   �  Ptype.func([]uint8, map[string]bool) bool   �  jtype.func(*"".Context, []uint8, map[string]bool) bool   �  2"".(*Context).shouldBuild   �  2"".(*Context).shouldBuild   �  :go.string.hdr."splitPathList"   �  "go.importpath."".   �  4type.func(string) []string   �  Ntype.func(*"".Context, string) []string   �  6"".(*Context).splitPathList   �  6"".(*Context).splitPathList   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[2]string              (type..hash.[2]string   �,type..eqfunc.[2]string              $type..eq.[2]string   �&type..alg.[2]string                        0type..hashfunc.[2]string     ,type..eqfunc.[2]string   �"runtime.gcbits.05    �2go.string.hdr."[2]string"             	          *go.string."[2]string"   �*go.string."[2]string"    [2]string  �type.[2]string �  �               PX��                                                                0  &type..alg.[2]string   @  "runtime.gcbits.05   P  2go.string.hdr."[2]string"   p  .go.weak.type.*[2]string   �  type.string   �  type.[]string   �>go.typelink.[2]string	[2]string              type.[2]string   �4go.string.hdr."*[2]string"             
          ,go.string."*[2]string"   �,go.string."*[2]string"    *[2]string  �type.*[2]string �  �              f< 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[2]string"   p  0go.weak.type.**[2]string   �  type.[2]string   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[6]string              (type..hash.[6]string   �,type..eqfunc.[6]string              $type..eq.[6]string   �&type..alg.[6]string                        0type..hashfunc.[6]string     ,type..eqfunc.[6]string   �&runtime.gcbits.5505   U �2go.string.hdr."[6]string"             	          *go.string."[6]string"   �*go.string."[6]string"    [6]string  �type.[6]string �  �`       X       �:�~                                                                0  &type..alg.[6]string   @  &runtime.gcbits.5505   P  2go.string.hdr."[6]string"   p  .go.weak.type.*[6]string   �  type.string   �  type.[]string   �>go.typelink.[6]string	[6]string              type.[6]string   �4go.string.hdr."*[6]string"             
          ,go.string."*[6]string"   �,go.string."*[6]string"    *[6]string  �type.*[6]string �  �              ��Y 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[6]string"   p  0go.weak.type.**[6]string   �  type.[6]string   � type..hashfunc32                        ,runtime.memhash_varlen   �type..eqfunc32                        .runtime.memequal_varlen   �type..alg32                         type..hashfunc32     type..eqfunc32   �2go.string.hdr."[32]uint8"             	          *go.string."[32]uint8"   �*go.string."[32]uint8"    [32]uint8  �type.[32]uint8 �  �                �Y�� �                                                                0  type..alg32   @  runtime.gcbits.   P  2go.string.hdr."[32]uint8"   p  .go.weak.type.*[32]uint8   �  type.uint8   �  type.[]uint8   �>go.typelink.[32]uint8	[32]uint8              type.[32]uint8   �>go.string.hdr."build.NoGoError"                       6go.string."build.NoGoError"   �6go.string."build.NoGoError"     build.NoGoError  �2go.string.hdr."NoGoError"             	          *go.string."NoGoError"   �*go.string."NoGoError"    NoGoError  �"type."".NoGoError  �  �              �s�@                                                                                                                                               0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."build.NoGoError"   p  $type.*"".NoGoError   �� "type."".NoGoError   �  &go.string.hdr."Dir"   �  type.string   `� "type."".NoGoError   �  2go.string.hdr."NoGoError"   �  "go.importpath."".   �� "type."".NoGoError   �@go.string.hdr."*build.NoGoError"                       8go.string."*build.NoGoError"   �8go.string."*build.NoGoError" 0  "*build.NoGoError  �Zgo.string.hdr."func(*build.NoGoError) string"                       Rgo.string."func(*build.NoGoError) string"   �Rgo.string."func(*build.NoGoError) string" @  <func(*build.NoGoError) string  �>type.func(*"".NoGoError) string �  �              �d� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."func(*build.NoGoError) string"   p  Pgo.weak.type.*func(*"".NoGoError) string   �� >type.func(*"".NoGoError) string   �� >type.func(*"".NoGoError) string   �  $type.*"".NoGoError   �  type.string   ��go.typelink.func(*build.NoGoError) string	func(*"".NoGoError) string              >type.func(*"".NoGoError) string   �*go.string.hdr."Error"                       "go.string."Error"   �"go.string."Error"   Error  �:go.string.hdr."func() string"                       2go.string."func() string"   �2go.string."func() string"    func() string  �$type.func() string �  �              �m� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."func() string"   p  6go.weak.type.*func() string   �� $type.func() string   �� $type.func() string   �  type.string   �Ngo.typelink.func() string	func() string              $type.func() string   �$type.*"".NoGoError  �  �              J�� 6                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*build.NoGoError"   p  6go.weak.type.**"".NoGoError   �  "type."".NoGoError   `� $type.*"".NoGoError   �� $type.*"".NoGoError   �  *go.string.hdr."Error"   �  $type.func() string   �  >type.func(*"".NoGoError) string   �  *"".(*NoGoError).Error   �  *"".(*NoGoError).Error   �"runtime.gcbits.25   % �Tgo.string.hdr."build.MultiplePackageError"                       Lgo.string."build.MultiplePackageError"   �Lgo.string."build.MultiplePackageError" @  6build.MultiplePackageError  �0go.string.hdr."Packages"                       (go.string."Packages"   �(go.string."Packages"    Packages  �*go.string.hdr."Files"                       "go.string."Files"   �"go.string."Files"   Files  �Hgo.string.hdr."MultiplePackageError"                       @go.string."MultiplePackageError"   �@go.string."MultiplePackageError" 0  *MultiplePackageError  �8type."".MultiplePackageError  �  �@       0       �27�                                                                                                                                                                              (                                               0�  runtime.algarray   @  "runtime.gcbits.25   P  Tgo.string.hdr."build.MultiplePackageError"   p  :type.*"".MultiplePackageError   �� 8type."".MultiplePackageError   �  &go.string.hdr."Dir"   �  type.string   �  0go.string.hdr."Packages"   �  type.[]string   �  *go.string.hdr."Files"   �  type.[]string   `� 8type."".MultiplePackageError   �  Hgo.string.hdr."MultiplePackageError"   �  "go.importpath."".   �� 8type."".MultiplePackageError   �Vgo.string.hdr."*build.MultiplePackageError"                       Ngo.string."*build.MultiplePackageError"   �Ngo.string."*build.MultiplePackageError" @  8*build.MultiplePackageError  �pgo.string.hdr."func(*build.MultiplePackageError) string"             (          hgo.string."func(*build.MultiplePackageError) string"   �hgo.string."func(*build.MultiplePackageError) string" `  Rfunc(*build.MultiplePackageError) string  �Ttype.func(*"".MultiplePackageError) string �  �              HM�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  pgo.string.hdr."func(*build.MultiplePackageError) string"   p  fgo.weak.type.*func(*"".MultiplePackageError) string   �� Ttype.func(*"".MultiplePackageError) string   �� Ttype.func(*"".MultiplePackageError) string   �  :type.*"".MultiplePackageError   �  type.string   ��go.typelink.func(*build.MultiplePackageError) string	func(*"".MultiplePackageError) string              Ttype.func(*"".MultiplePackageError) string   �:type.*"".MultiplePackageError  �  �              o�R� 6                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Vgo.string.hdr."*build.MultiplePackageError"   p  Lgo.weak.type.**"".MultiplePackageError   �  8type."".MultiplePackageError   `� :type.*"".MultiplePackageError   �� :type.*"".MultiplePackageError   �  *go.string.hdr."Error"   �  $type.func() string   �  Ttype.func(*"".MultiplePackageError) string   �  @"".(*MultiplePackageError).Error   �  @"".(*MultiplePackageError).Error   �"runtime.gcbits.03    �8go.string.hdr."interface {}"                       0go.string."interface {}"   �0go.string."interface {}"    interface {}  �"type.interface {} �  �              �W�                                                                 
0�  runtime.algarray   @  "runtime.gcbits.03   P  8go.string.hdr."interface {}"   p  4go.weak.type.*interface {}   �� "type.interface {}   �<go.string.hdr."[]interface {}"                       4go.string."[]interface {}"   �4go.string."[]interface {}"    []interface {}  �&type.[]interface {} �  �              p��/                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."[]interface {}"   p  8go.weak.type.*[]interface {}   �  "type.interface {}   �Rgo.typelink.[]interface {}	[]interface {}              &type.[]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[5]interface {}              4type..hash.[5]interface {}   �8type..eqfunc.[5]interface {}              0type..eq.[5]interface {}   �2type..alg.[5]interface {}                        <type..hashfunc.[5]interface {}     8type..eqfunc.[5]interface {}   �&runtime.gcbits.ff03   � �>go.string.hdr."[5]interface {}"                       6go.string."[5]interface {}"   �6go.string."[5]interface {}"     [5]interface {}  �(type.[5]interface {} �  �P       P       �#��                                                                0  2type..alg.[5]interface {}   @  &runtime.gcbits.ff03   P  >go.string.hdr."[5]interface {}"   p  :go.weak.type.*[5]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[5]interface {}	[5]interface {}              (type.[5]interface {}   �@go.string.hdr."*[5]interface {}"                       8go.string."*[5]interface {}"   �8go.string."*[5]interface {}" 0  "*[5]interface {}  �*type.*[5]interface {} �  �              �?@ 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[5]interface {}"   p  <go.weak.type.**[5]interface {}   �  (type.[5]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[3]string              (type..hash.[3]string   �,type..eqfunc.[3]string              $type..eq.[3]string   �&type..alg.[3]string                        0type..hashfunc.[3]string     ,type..eqfunc.[3]string   �"runtime.gcbits.15    �2go.string.hdr."[3]string"             	          *go.string."[3]string"   �*go.string."[3]string"    [3]string  �type.[3]string �  �0       (       C�iB                                                                0  &type..alg.[3]string   @  "runtime.gcbits.15   P  2go.string.hdr."[3]string"   p  .go.weak.type.*[3]string   �  type.string   �  type.[]string   �>go.typelink.[3]string	[3]string              type.[3]string   �,go.string.hdr."func()"                       $go.string."func()"   �$go.string."func()"   func()  �type.func() �  �              ���� 3                                                                                                0�  runtime.algarray   @  "runtime.gcbits.01   P  ,go.string.hdr."func()"   p  (go.weak.type.*func()   �� type.func()   �� type.func()   �2go.typelink.func()	func()              type.func()   �"runtime.gcbits.29   ) ��go.string.hdr."struct { vendor []string; goroot string; gopath []string }"             :          �go.string."struct { vendor []string; goroot string; gopath []string }"   ��go.string."struct { vendor []string; goroot string; gopath []string }" �  vstruct { vendor []string; goroot string; gopath []string }  �,go.string.hdr."goroot"                       $go.string."goroot"   �$go.string."goroot"   goroot  �~type.struct { vendor []string; goroot string; gopath []string } �  �@       0       �q�D                                                                                                                                                                              (       0�  runtime.algarray   @  "runtime.gcbits.29   P  �go.string.hdr."struct { vendor []string; goroot string; gopath []string }"   p  �go.weak.type.*struct { vendor []string; goroot string; gopath []string }   �� ~type.struct { vendor []string; goroot string; gopath []string }   �  ,go.string.hdr."vendor"   �  "go.importpath."".   �  type.[]string   �  ,go.string.hdr."goroot"   �  "go.importpath."".   �  type.string   �  ,go.string.hdr."gopath"   �  "go.importpath."".   �  type.[]string   �Ngo.string.hdr."func(string, bool) bool"                       Fgo.string."func(string, bool) bool"   �Fgo.string."func(string, bool) bool" 0  0func(string, bool) bool  �8type.func(string, bool) bool �  �              g*n� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."func(string, bool) bool"   p  Jgo.weak.type.*func(string, bool) bool   �� 8type.func(string, bool) bool   �� 8type.func(string, bool) bool   �  type.string   �  type.bool   �  type.bool   �vgo.typelink.func(string, bool) bool	func(string, bool) bool              8type.func(string, bool) bool   �6go.string.hdr."func(error)"                       .go.string."func(error)"   �.go.string."func(error)"    func(error)  � type.func(error) �  �              ['g 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."func(error)"   p  2go.weak.type.*func(error)   ��  type.func(error)   ��  type.func(error)   �  type.error   �Fgo.typelink.func(error)	func(error)               type.func(error)   �4go.string.hdr."[]ast.Decl"             
          ,go.string."[]ast.Decl"   �,go.string."[]ast.Decl"    []ast.Decl  �$type.[]go/ast.Decl �  �              q|�+                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."[]ast.Decl"   p  6go.weak.type.*[]go/ast.Decl   �   type.go/ast.Decl   �Hgo.typelink.[]ast.Decl	[]go/ast.Decl              $type.[]go/ast.Decl   �4go.string.hdr."[]ast.Spec"             
          ,go.string."[]ast.Spec"   �,go.string."[]ast.Spec"    []ast.Spec  �$type.[]go/ast.Spec �  �              0�4                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."[]ast.Spec"   p  6go.weak.type.*[]go/ast.Spec   �   type.go/ast.Spec   �Hgo.typelink.[]ast.Spec	[]go/ast.Spec              $type.[]go/ast.Spec   �Hgo.string.hdr."*map.hdr[string]bool"                       @go.string."*map.hdr[string]bool"   �@go.string."*map.hdr[string]bool" 0  **map.hdr[string]bool  �2type.*map.hdr[string]bool �  �              ~� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."*map.hdr[string]bool"   p  Dgo.weak.type.**map.hdr[string]bool   �  0type.map.hdr[string]bool   �"runtime.gcbits.ff   � �Hgo.string.hdr."map.iter[string]bool"                       @go.string."map.iter[string]bool"   �@go.string."map.iter[string]bool" 0  *map.iter[string]bool  �&go.string.hdr."key"                       go.string."key"   �go.string."key"   key  �&go.string.hdr."val"                       go.string."val"   �go.string."val"   val  �"go.string.hdr."t"                       go.string."t"   �go.string."t"   t  �"go.string.hdr."h"                       go.string."h"   �go.string."h"   h  �(go.string.hdr."bptr"                        go.string."bptr"   � go.string."bptr"   
bptr  �2go.string.hdr."overflow0"             	          *go.string."overflow0"   �*go.string."overflow0"    overflow0  �2go.string.hdr."overflow1"             	          *go.string."overflow1"   �*go.string."overflow1"    overflow1  �6go.string.hdr."startBucket"                       .go.string."startBucket"   �.go.string."startBucket"    startBucket  �*go.string.hdr."stuff"                       "go.string."stuff"   �"go.string."stuff"   stuff  �,go.string.hdr."bucket"                       $go.string."bucket"   �$go.string."bucket"   bucket  �6go.string.hdr."checkBucket"                       .go.string."checkBucket"   �.go.string."checkBucket"    checkBucket  �2type.map.iter[string]bool �  �`       @       Q���                                                                                                                                                                                                                                                                                                    (                                       0                                       8                                       @                                       H                                       P                                       X       :0�  runtime.algarray   @  "runtime.gcbits.ff   P  Hgo.string.hdr."map.iter[string]bool"   p  Dgo.weak.type.*map.iter[string]bool   �� 2type.map.iter[string]bool   �  &go.string.hdr."key"   �  type.*string   �  &go.string.hdr."val"   �  type.*bool   �  "go.string.hdr."t"   �  type.*uint8   �  "go.string.hdr."h"   �  2type.*map.hdr[string]bool   �  .go.string.hdr."buckets"   �  8type.*map.bucket[string]bool   �  (go.string.hdr."bptr"   �  8type.*map.bucket[string]bool   �  2go.string.hdr."overflow0"   �  &type.unsafe.Pointer   �  2go.string.hdr."overflow1"   �  &type.unsafe.Pointer   �  6go.string.hdr."startBucket"   �  type.uintptr   �  *go.string.hdr."stuff"   �  type.uintptr   �  ,go.string.hdr."bucket"   �  type.uintptr   �  6go.string.hdr."checkBucket"   �  type.uintptr   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[1]interface {}              4type..hash.[1]interface {}   �8type..eqfunc.[1]interface {}              0type..eq.[1]interface {}   �2type..alg.[1]interface {}                        <type..hashfunc.[1]interface {}     8type..eqfunc.[1]interface {}   �>go.string.hdr."[1]interface {}"                       6go.string."[1]interface {}"   �6go.string."[1]interface {}"     [1]interface {}  �(type.[1]interface {} �  �              P�[�                                                                0  2type..alg.[1]interface {}   @  "runtime.gcbits.03   P  >go.string.hdr."[1]interface {}"   p  :go.weak.type.*[1]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[1]interface {}	[1]interface {}              (type.[1]interface {}   �@go.string.hdr."*[1]interface {}"                       8go.string."*[1]interface {}"   �8go.string."*[1]interface {}" 0  "*[1]interface {}  �*type.*[1]interface {} �  �              ��5 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[1]interface {}"   p  <go.weak.type.**[1]interface {}   �  (type.[1]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[2]interface {}              4type..hash.[2]interface {}   �8type..eqfunc.[2]interface {}              0type..eq.[2]interface {}   �2type..alg.[2]interface {}                        <type..hashfunc.[2]interface {}     8type..eqfunc.[2]interface {}   �"runtime.gcbits.0f    �>go.string.hdr."[2]interface {}"                       6go.string."[2]interface {}"   �6go.string."[2]interface {}"     [2]interface {}  �(type.[2]interface {} �  �                ,Y��                                                                0  2type..alg.[2]interface {}   @  "runtime.gcbits.0f   P  >go.string.hdr."[2]interface {}"   p  :go.weak.type.*[2]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[2]interface {}	[2]interface {}              (type.[2]interface {}   �@go.string.hdr."*[2]interface {}"                       8go.string."*[2]interface {}"   �8go.string."*[2]interface {}" 0  "*[2]interface {}  �*type.*[2]interface {} �  �              �s-q 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[2]interface {}"   p  <go.weak.type.**[2]interface {}   �  (type.[2]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             ��type..hashfunc.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }              �type..hash.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   ��type..eqfunc.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }              �type..eq.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   ��type..alg.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }                        �type..hashfunc.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }     �type..eqfunc.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   �"runtime.gcbits.1e    ��go.string.hdr."struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"             _          �go.string."struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"   ��go.string."struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }" �  �struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }  �$go.string.hdr.".F"                       go.string.".F"   �go.string.".F"   .F  �(go.string.hdr."ctxt"                        go.string."ctxt"   � go.string."ctxt"   
ctxt  �"go.string.hdr."p"                       go.string."p"   �go.string."p"   p  �(go.string.hdr."pkga"                        go.string."pkga"   � go.string."pkga"   
pkga  �:go.string.hdr."pkgtargetroot"                       2go.string."pkgtargetroot"   �2go.string."pkgtargetroot"    pkgtargetroot  ��type.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } �  �0       (       x<K}                                                                                                                                                                                                                                                                    (0  �type..alg.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   @  "runtime.gcbits.1e   P  �go.string.hdr."struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"   p  �go.weak.type.*struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   �� �type.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   �  $go.string.hdr.".F"   �  "go.importpath."".   �  type.uintptr   �  (go.string.hdr."ctxt"   �  "go.importpath."".   �   type.*"".Context   �  "go.string.hdr."p"   �  "go.importpath."".   �   type.*"".Package   �  (go.string.hdr."pkga"   �  "go.importpath."".   �  type.*string   �  :go.string.hdr."pkgtargetroot"   �  "go.importpath."".   �  type.string   ��go.string.hdr."*struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"             `          �go.string."*struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"   ��go.string."*struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }" �  �*struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }  ��type.*struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string } �  �              P�a� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."*struct { F uintptr; ctxt *build.Context; p *build.Package; pkga *string; pkgtargetroot string }"   p  �go.weak.type.**struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   �  �type.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   �4go.string.hdr."*[3]string"             
          ,go.string."*[3]string"   �,go.string."*[3]string"    *[3]string  �type.*[3]string �  �              
+� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[3]string"   p  0go.weak.type.**[3]string   �  type.[3]string   ��go.string.hdr."*struct { vendor []string; goroot string; gopath []string }"             ;          �go.string."*struct { vendor []string; goroot string; gopath []string }"   ��go.string."*struct { vendor []string; goroot string; gopath []string }" �  x*struct { vendor []string; goroot string; gopath []string }  ��type.*struct { vendor []string; goroot string; gopath []string } �  �              ��% 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."*struct { vendor []string; goroot string; gopath []string }"   p  �go.weak.type.**struct { vendor []string; goroot string; gopath []string }   �  ~type.struct { vendor []string; goroot string; gopath []string }   �&runtime.gcbits.d601   � �$"".hdr..gostring.2             �          ""..gostring.2   �""..gostring.2 �  �struct { F uintptr; ctxt *build.Context; srcDir string; path string; p *build.Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }  �,go.string.hdr."srcDir"                       $go.string."srcDir"   �$go.string."srcDir"   srcDir  �(go.string.hdr."path"                        go.string."path"   � go.string."path"   
path  �.go.string.hdr."setPkga"                       &go.string."setPkga"   �&go.string."setPkga"   setPkga  �*go.string.hdr."tried"                       "go.string."tried"   �"go.string."tried"   tried  ��type.struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } } �  �H       H       *e��                                                                                                                                                                                                                                                             0                                       8                                       @       40�  runtime.algarray   @  &runtime.gcbits.d601   P  $"".hdr..gostring.2   p  �go.weak.type.*struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }   �� �type.struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }   �  $go.string.hdr.".F"   �  "go.importpath."".   �  type.uintptr   �  (go.string.hdr."ctxt"   �  "go.importpath."".   �   type.*"".Context   �  ,go.string.hdr."srcDir"   �  "go.importpath."".   �  type.string   �  (go.string.hdr."path"   �  "go.importpath."".   �  type.string   �  "go.string.hdr."p"   �  "go.importpath."".   �   type.*"".Package   �  .go.string.hdr."setPkga"   �  "go.importpath."".   �  type.func()   �  *go.string.hdr."tried"   �  "go.importpath."".   �  �type.*struct { vendor []string; goroot string; gopath []string }   �$"".hdr..gostring.3             �          ""..gostring.3   �""..gostring.3 �  �*struct { F uintptr; ctxt *build.Context; srcDir string; path string; p *build.Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }  ��type.*struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } } �  �              �v 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  $"".hdr..gostring.3   p  �go.weak.type.**struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }   �  �type.struct { F uintptr; ctxt *"".Context; srcDir string; path string; p *"".Package; setPkga func(); tried *struct { vendor []string; goroot string; gopath []string } }   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             ��type..hashfunc.struct { F uintptr; badGoError *error; p *"".Package; name string }              �type..hash.struct { F uintptr; badGoError *error; p *"".Package; name string }   ��type..eqfunc.struct { F uintptr; badGoError *error; p *"".Package; name string }              �type..eq.struct { F uintptr; badGoError *error; p *"".Package; name string }   ��type..alg.struct { F uintptr; badGoError *error; p *"".Package; name string }                        �type..hashfunc.struct { F uintptr; badGoError *error; p *"".Package; name string }     �type..eqfunc.struct { F uintptr; badGoError *error; p *"".Package; name string }   �"runtime.gcbits.0e    ��go.string.hdr."struct { F uintptr; badGoError *error; p *build.Package; name string }"             F          �go.string."struct { F uintptr; badGoError *error; p *build.Package; name string }"   ��go.string."struct { F uintptr; badGoError *error; p *build.Package; name string }" �  �struct { F uintptr; badGoError *error; p *build.Package; name string }  �4go.string.hdr."badGoError"             
          ,go.string."badGoError"   �,go.string."badGoError"    badGoError  �(go.string.hdr."name"                        go.string."name"   � go.string."name"   
name  ��type.struct { F uintptr; badGoError *error; p *"".Package; name string } �  �(               ��JE                                                                                                                                                                                                                            "0  �type..alg.struct { F uintptr; badGoError *error; p *"".Package; name string }   @  "runtime.gcbits.0e   P  �go.string.hdr."struct { F uintptr; badGoError *error; p *build.Package; name string }"   p  �go.weak.type.*struct { F uintptr; badGoError *error; p *"".Package; name string }   �� �type.struct { F uintptr; badGoError *error; p *"".Package; name string }   �  $go.string.hdr.".F"   �  "go.importpath."".   �  type.uintptr   �  4go.string.hdr."badGoError"   �  "go.importpath."".   �  type.*error   �  "go.string.hdr."p"   �  "go.importpath."".   �   type.*"".Package   �  (go.string.hdr."name"   �  "go.importpath."".   �  type.string   ��go.string.hdr."*struct { F uintptr; badGoError *error; p *build.Package; name string }"             G          �go.string."*struct { F uintptr; badGoError *error; p *build.Package; name string }"   ��go.string."*struct { F uintptr; badGoError *error; p *build.Package; name string }" �  �*struct { F uintptr; badGoError *error; p *build.Package; name string }  ��type.*struct { F uintptr; badGoError *error; p *"".Package; name string } �  �              m�� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."*struct { F uintptr; badGoError *error; p *build.Package; name string }"   p  �go.weak.type.**struct { F uintptr; badGoError *error; p *"".Package; name string }   �  �type.struct { F uintptr; badGoError *error; p *"".Package; name string }   �Bgo.string.hdr."*[]token.Position"                       :go.string."*[]token.Position"   �:go.string."*[]token.Position" 0  $*[]token.Position  �2type.*[]go/token.Position �  �              ^+� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."*[]token.Position"   p  Dgo.weak.type.**[]go/token.Position   �  0type.[]go/token.Position   �`go.string.hdr."*map.hdr[string][]token.Position"                        Xgo.string."*map.hdr[string][]token.Position"   �Xgo.string."*map.hdr[string][]token.Position" P  B*map.hdr[string][]token.Position  �Ptype.*map.hdr[string][]go/token.Position �  �              �u� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."*map.hdr[string][]token.Position"   p  bgo.weak.type.**map.hdr[string][]go/token.Position   �  Ntype.map.hdr[string][]go/token.Position   �`go.string.hdr."map.iter[string][]token.Position"                        Xgo.string."map.iter[string][]token.Position"   �Xgo.string."map.iter[string][]token.Position" P  Bmap.iter[string][]token.Position  �Ptype.map.iter[string][]go/token.Position �  �`       @       .���                                                                                                                                                                                                                                                                                                    (                                       0                                       8                                       @                                       H                                       P                                       X       :0�  runtime.algarray   @  "runtime.gcbits.ff   P  `go.string.hdr."map.iter[string][]token.Position"   p  bgo.weak.type.*map.iter[string][]go/token.Position   �� Ptype.map.iter[string][]go/token.Position   �  &go.string.hdr."key"   �  type.*string   �  &go.string.hdr."val"   �  2type.*[]go/token.Position   �  "go.string.hdr."t"   �  type.*uint8   �  "go.string.hdr."h"   �  Ptype.*map.hdr[string][]go/token.Position   �  .go.string.hdr."buckets"   �  Vtype.*map.bucket[string][]go/token.Position   �  (go.string.hdr."bptr"   �  Vtype.*map.bucket[string][]go/token.Position   �  2go.string.hdr."overflow0"   �  &type.unsafe.Pointer   �  2go.string.hdr."overflow1"   �  &type.unsafe.Pointer   �  6go.string.hdr."startBucket"   �  type.uintptr   �  *go.string.hdr."stuff"   �  type.uintptr   �  ,go.string.hdr."bucket"   �  type.uintptr   �  6go.string.hdr."checkBucket"   �  type.uintptr   �.go.string.hdr."[]int32"                       &go.string."[]int32"   �&go.string."[]int32"   []int32  �type.[]int32 �  �              *Ms                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  .go.string.hdr."[]int32"   p  *go.weak.type.*[]int32   �  type.int32   �6go.typelink.[]int32	[]int32              type.[]int32   �"runtime.gcbits.63   c �Dgo.string.hdr."build.importReader"                       <go.string."build.importReader"   �<go.string."build.importReader" 0  &build.importReader  �"go.string.hdr."b"                       go.string."b"   �go.string."b"   b  �&go.string.hdr."buf"                       go.string."buf"   �go.string."buf"   buf  �(go.string.hdr."peek"                        go.string."peek"   � go.string."peek"   
peek  �&go.string.hdr."err"                       go.string."err"   �go.string."err"   err  �&go.string.hdr."eof"                       go.string."eof"   �go.string."eof"   eof  �(go.string.hdr."nerr"                        go.string."nerr"   � go.string."nerr"   
nerr  �8go.string.hdr."importReader"                       0go.string."importReader"   �0go.string."importReader"    importReader  �(type."".importReader  �  �H       8       �K}a                                                                                                                                                                                                                      (                                       8                                       @                                               60�  runtime.algarray   @  "runtime.gcbits.63   P  Dgo.string.hdr."build.importReader"   p  *type.*"".importReader   �� (type."".importReader   �  "go.string.hdr."b"   �  "go.importpath."".   �  $type.*bufio.Reader   �  &go.string.hdr."buf"   �  "go.importpath."".   �  type.[]uint8   �  (go.string.hdr."peek"   �  "go.importpath."".   �  type.uint8   �  &go.string.hdr."err"   �  "go.importpath."".   �  type.error   �  &go.string.hdr."eof"   �  "go.importpath."".   �  type.bool   �  (go.string.hdr."nerr"   �  "go.importpath."".   �  type.int   `� (type."".importReader   �  8go.string.hdr."importReader"   �  "go.importpath."".   �� (type."".importReader   �Fgo.string.hdr."*build.importReader"                       >go.string."*build.importReader"   �>go.string."*build.importReader" 0  (*build.importReader  �jgo.string.hdr."func(*build.importReader, bool) uint8"             %          bgo.string."func(*build.importReader, bool) uint8"   �bgo.string."func(*build.importReader, bool) uint8" P  Lfunc(*build.importReader, bool) uint8  �Ntype.func(*"".importReader, bool) uint8 �  �              F�� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(*build.importReader, bool) uint8"   p  `go.weak.type.*func(*"".importReader, bool) uint8   �� Ntype.func(*"".importReader, bool) uint8   �� Ntype.func(*"".importReader, bool) uint8   �  *type.*"".importReader   �  type.bool   �  type.uint8   ��go.typelink.func(*build.importReader, bool) uint8	func(*"".importReader, bool) uint8              Ntype.func(*"".importReader, bool) uint8   �^go.string.hdr."func(*build.importReader) uint8"                       Vgo.string."func(*build.importReader) uint8"   �Vgo.string."func(*build.importReader) uint8" @  @func(*build.importReader) uint8  �Btype.func(*"".importReader) uint8 �  �              _�2 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(*build.importReader) uint8"   p  Tgo.weak.type.*func(*"".importReader) uint8   �� Btype.func(*"".importReader) uint8   �� Btype.func(*"".importReader) uint8   �  *type.*"".importReader   �  type.uint8   ��go.typelink.func(*build.importReader) uint8	func(*"".importReader) uint8              Btype.func(*"".importReader) uint8   �Rgo.string.hdr."func(*build.importReader)"                       Jgo.string."func(*build.importReader)"   �Jgo.string."func(*build.importReader)" @  4func(*build.importReader)  �6type.func(*"".importReader) �  �              5�;& 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func(*build.importReader)"   p  Hgo.weak.type.*func(*"".importReader)   �� 6type.func(*"".importReader)   �� 6type.func(*"".importReader)   �  *type.*"".importReader   �xgo.typelink.func(*build.importReader)	func(*"".importReader)              6type.func(*"".importReader)   �2go.string.hdr."*[]string"             	          *go.string."*[]string"   �*go.string."*[]string"    *[]string  �type.*[]string �  �              �"v� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*[]string"   p  .go.weak.type.**[]string   �  type.[]string   �hgo.string.hdr."func(*build.importReader, *[]string)"             $          `go.string."func(*build.importReader, *[]string)"   �`go.string."func(*build.importReader, *[]string)" P  Jfunc(*build.importReader, *[]string)  �Ltype.func(*"".importReader, *[]string) �  �              �ib 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  hgo.string.hdr."func(*build.importReader, *[]string)"   p  ^go.weak.type.*func(*"".importReader, *[]string)   �� Ltype.func(*"".importReader, *[]string)   �� Ltype.func(*"".importReader, *[]string)   �  *type.*"".importReader   �  type.*[]string   ��go.typelink.func(*build.importReader, *[]string)	func(*"".importReader, *[]string)              Ltype.func(*"".importReader, *[]string)   �bgo.string.hdr."func(*build.importReader, string)"             !          Zgo.string."func(*build.importReader, string)"   �Zgo.string."func(*build.importReader, string)" P  Dfunc(*build.importReader, string)  �Ftype.func(*"".importReader, string) �  �              `�|� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*build.importReader, string)"   p  Xgo.weak.type.*func(*"".importReader, string)   �� Ftype.func(*"".importReader, string)   �� Ftype.func(*"".importReader, string)   �  *type.*"".importReader   �  type.string   ��go.typelink.func(*build.importReader, string)	func(*"".importReader, string)              Ftype.func(*"".importReader, string)   �0go.string.hdr."nextByte"                       (go.string."nextByte"   �(go.string."nextByte"    nextByte  �@go.string.hdr."func(bool) uint8"                       8go.string."func(bool) uint8"   �8go.string."func(bool) uint8" 0  "func(bool) uint8  �*type.func(bool) uint8 �  �              �j� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."func(bool) uint8"   p  <go.weak.type.*func(bool) uint8   �� *type.func(bool) uint8   �� *type.func(bool) uint8   �  type.bool   �  type.uint8   �Zgo.typelink.func(bool) uint8	func(bool) uint8              *type.func(bool) uint8   �0go.string.hdr."peekByte"                       (go.string."peekByte"   �(go.string."peekByte"    peekByte  �0go.string.hdr."readByte"                       (go.string."readByte"   �(go.string."readByte"    readByte  �8go.string.hdr."func() uint8"                       0go.string."func() uint8"   �0go.string."func() uint8"    func() uint8  �"type.func() uint8 �  �              }S'� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."func() uint8"   p  4go.weak.type.*func() uint8   �� "type.func() uint8   �� "type.func() uint8   �  type.uint8   �Jgo.typelink.func() uint8	func() uint8              "type.func() uint8   �2go.string.hdr."readIdent"             	          *go.string."readIdent"   �*go.string."readIdent"    readIdent  �4go.string.hdr."readImport"             
          ,go.string."readImport"   �,go.string."readImport"    readImport  �>go.string.hdr."func(*[]string)"                       6go.string."func(*[]string)"   �6go.string."func(*[]string)"     func(*[]string)  �(type.func(*[]string) �  �              �ު 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."func(*[]string)"   p  :go.weak.type.*func(*[]string)   �� (type.func(*[]string)   �� (type.func(*[]string)   �  type.*[]string   �Vgo.typelink.func(*[]string)	func(*[]string)              (type.func(*[]string)   �6go.string.hdr."readKeyword"                       .go.string."readKeyword"   �.go.string."readKeyword"    readKeyword  �8go.string.hdr."func(string)"                       0go.string."func(string)"   �0go.string."func(string)"    func(string)  �"type.func(string) �  �              �ǹ� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."func(string)"   p  4go.weak.type.*func(string)   �� "type.func(string)   �� "type.func(string)   �  type.string   �Jgo.typelink.func(string)	func(string)              "type.func(string)   �4go.string.hdr."readString"             
          ,go.string."readString"   �,go.string."readString"    readString  �6go.string.hdr."syntaxError"                       .go.string."syntaxError"   �.go.string."syntaxError"    syntaxError  �*type.*"".importReader  �  �              �p�� 6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      n0�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."*build.importReader"   p  <go.weak.type.**"".importReader   �  (type."".importReader   `� *type.*"".importReader   �� *type.*"".importReader   �  0go.string.hdr."nextByte"   �  "go.importpath."".   �  *type.func(bool) uint8   �  Ntype.func(*"".importReader, bool) uint8   �  6"".(*importReader).nextByte   �  6"".(*importReader).nextByte   �  0go.string.hdr."peekByte"   �  "go.importpath."".   �  *type.func(bool) uint8   �  Ntype.func(*"".importReader, bool) uint8   �  6"".(*importReader).peekByte   �  6"".(*importReader).peekByte   �  0go.string.hdr."readByte"   �  "go.importpath."".   �  "type.func() uint8   �  Btype.func(*"".importReader) uint8   �  6"".(*importReader).readByte   �  6"".(*importReader).readByte   �  2go.string.hdr."readIdent"   �  "go.importpath."".   �  type.func()   �  6type.func(*"".importReader)   �  8"".(*importReader).readIdent   �  8"".(*importReader).readIdent   �  4go.string.hdr."readImport"   �  "go.importpath."".   �  (type.func(*[]string)   �  Ltype.func(*"".importReader, *[]string)   �  :"".(*importReader).readImport   �  :"".(*importReader).readImport   �  6go.string.hdr."readKeyword"   �  "go.importpath."".   �  "type.func(string)   �  Ftype.func(*"".importReader, string)   �  <"".(*importReader).readKeyword   �  <"".(*importReader).readKeyword   �  4go.string.hdr."readString"   �  "go.importpath."".   �  (type.func(*[]string)   �  Ltype.func(*"".importReader, *[]string)   �  :"".(*importReader).readString   �  :"".(*importReader).readString   �  6go.string.hdr."syntaxError"   �  "go.importpath."".   �  type.func()   �  6type.func(*"".importReader)   �  <"".(*importReader).syntaxError   �  <"".(*importReader).syntaxError   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �Ttype..hashfunc.struct { a string; b bool }              Ltype..hash.struct { a string; b bool }   �Ptype..eqfunc.struct { a string; b bool }              Htype..eq.struct { a string; b bool }   �Jtype..alg.struct { a string; b bool }                        Ttype..hashfunc.struct { a string; b bool }     Ptype..eqfunc.struct { a string; b bool }   �Vgo.string.hdr."struct { a string; b bool }"                       Ngo.string."struct { a string; b bool }"   �Ngo.string."struct { a string; b bool }" @  8struct { a string; b bool }  �"go.string.hdr."a"                       go.string."a"   �go.string."a"   a  �@type.struct { a string; b bool } �  �              ��                                                                                                                                              0  Jtype..alg.struct { a string; b bool }   @  "runtime.gcbits.01   P  Vgo.string.hdr."struct { a string; b bool }"   p  Rgo.weak.type.*struct { a string; b bool }   �� @type.struct { a string; b bool }   �  "go.string.hdr."a"   �  "go.importpath."".   �  type.string   �  "go.string.hdr."b"   �  "go.importpath."".   �  type.bool   �Zgo.string.hdr."[]struct { a string; b bool }"                       Rgo.string."[]struct { a string; b bool }"   �Rgo.string."[]struct { a string; b bool }" @  <[]struct { a string; b bool }  �Dtype.[]struct { a string; b bool } �  �              ��M�                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."[]struct { a string; b bool }"   p  Vgo.weak.type.*[]struct { a string; b bool }   �  @type.struct { a string; b bool }   ��go.typelink.[]struct { a string; b bool }	[]struct { a string; b bool }              Dtype.[]struct { a string; b bool }   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·34eab47d33fa46b254c22cdccfd2dc77                   �Tgclocals·51af24152615272c3d9efc8538f95767                  �\type..hashfunc.[24]struct { a string; b bool }              Ttype..hash.[24]struct { a string; b bool }   �Xtype..eqfunc.[24]struct { a string; b bool }              Ptype..eq.[24]struct { a string; b bool }   �Rtype..alg.[24]struct { a string; b bool }                        \type..hashfunc.[24]struct { a string; b bool }     Xtype..eqfunc.[24]struct { a string; b bool }   �Bruntime.gcbits.499224499224499224   I�$I�$I�$ �^go.string.hdr."[24]struct { a string; b bool }"                       Vgo.string."[24]struct { a string; b bool }"   �Vgo.string."[24]struct { a string; b bool }" @  @[24]struct { a string; b bool }  �Htype.[24]struct { a string; b bool } �  �@      0      �P��                                                                0  Rtype..alg.[24]struct { a string; b bool }   @  Bruntime.gcbits.499224499224499224   P  ^go.string.hdr."[24]struct { a string; b bool }"   p  Zgo.weak.type.*[24]struct { a string; b bool }   �  @type.struct { a string; b bool }   �  Dtype.[]struct { a string; b bool }   ��go.typelink.[24]struct { a string; b bool }	[24]struct { a string; b bool }              Htype.[24]struct { a string; b bool }   �4go.string.hdr."*[8]string"             
          ,go.string."*[8]string"   �,go.string."*[8]string"    *[8]string  �type.*[8]string �  �              ��o 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[8]string"   p  0go.weak.type.**[8]string   �  type.[8]string   �Xgo.string.hdr."*struct { a string; b bool }"                       Pgo.string."*struct { a string; b bool }"   �Pgo.string."*struct { a string; b bool }" @  :*struct { a string; b bool }  �Btype.*struct { a string; b bool } �  �              �c� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."*struct { a string; b bool }"   p  Tgo.weak.type.**struct { a string; b bool }   �  @type.struct { a string; b bool }   �`go.string.hdr."*[24]struct { a string; b bool }"                        Xgo.string."*[24]struct { a string; b bool }"   �Xgo.string."*[24]struct { a string; b bool }" P  B*[24]struct { a string; b bool }  �Jtype.*[24]struct { a string; b bool } �  �              ߷� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."*[24]struct { a string; b bool }"   p  \go.weak.type.**[24]struct { a string; b bool }   �  Htype.[24]struct { a string; b bool }   �.go.string.hdr."runtime"                       &go.string."runtime"   �&go.string."runtime"   runtime  �,go.importpath.runtime.                       &go.string."runtime"   �*go.string.hdr."bytes"                       "go.string."bytes"   �"go.string."bytes"   bytes  �(go.importpath.bytes.                       "go.string."bytes"   �,go.string.hdr."errors"                       $go.string."errors"   �$go.string."errors"   errors  �*go.importpath.errors.                       $go.string."errors"   �$go.string.hdr."io"                       go.string."io"   �go.string."io"   io  �"go.importpath.io.                       go.string."io"   �8go.string.hdr."unicode/utf8"                       0go.string."unicode/utf8"   �0go.string."unicode/utf8"    unicode/utf8  �6go.importpath.unicode/utf8.                       0go.string."unicode/utf8"   �.go.string.hdr."unicode"                       &go.string."unicode"   �&go.string."unicode"   unicode  �,go.importpath.unicode.                       &go.string."unicode"   �&go.string.hdr."fmt"                       go.string."fmt"   �go.string."fmt"   fmt  �$go.importpath.fmt.                       go.string."fmt"   �.go.string.hdr."strconv"                       &go.string."strconv"   �&go.string."strconv"   strconv  �,go.importpath.strconv.                       &go.string."strconv"   �$go.string.hdr."os"                       go.string."os"   �go.string."os"   os  �"go.importpath.os.                       go.string."os"   �,go.string.hdr."go/ast"                       $go.string."go/ast"   �$go.string."go/ast"   go/ast  �*go.importpath.go/ast.                       $go.string."go/ast"   �0go.string.hdr."go/token"                       (go.string."go/token"   �(go.string."go/token"    go/token  �.go.importpath.go/token.                       (go.string."go/token"   �(go.string.hdr."sort"                        go.string."sort"   � go.string."sort"   
sort  �&go.importpath.sort.                        go.string."sort"   �.go.string.hdr."strings"                       &go.string."strings"   �&go.string."strings"   strings  �,go.importpath.strings.                       &go.string."strings"   �,go.string.hdr."go/doc"                       $go.string."go/doc"   �$go.string."go/doc"   go/doc  �*go.importpath.go/doc.                       $go.string."go/doc"   �&go.importpath.path.                        go.string."path"   �2go.string.hdr."go/parser"             	          *go.string."go/parser"   �*go.string."go/parser"    go/parser  �0go.importpath.go/parser.             	          *go.string."go/parser"   �2go.string.hdr."io/ioutil"             	          *go.string."io/ioutil"   �*go.string."io/ioutil"    io/ioutil  �0go.importpath.io/ioutil.             	          *go.string."io/ioutil"   �:go.string.hdr."path/filepath"                       2go.string."path/filepath"   �2go.string."path/filepath"    path/filepath  �8go.importpath.path/filepath.                       2go.string."path/filepath"   �&go.string.hdr."log"                       go.string."log"   �go.string."log"   log  �$go.importpath.log.                       go.string."log"   �*go.string.hdr."bufio"                       "go.string."bufio"   �"go.string."bufio"   bufio  �(go.importpath.bufio.                       "go.string."bufio"   �.type..hash.[8]string·f              (type..hash.[8]string   �*type..eq.[8]string·f              $type..eq.[8]string   �.type..hash.[2]string·f              (type..hash.[2]string   �*type..eq.[2]string·f              $type..eq.[2]string   �.type..hash.[6]string·f              (type..hash.[6]string   �*type..eq.[6]string·f              $type..eq.[6]string   �:type..hash.[5]interface {}·f              4type..hash.[5]interface {}   �6type..eq.[5]interface {}·f              0type..eq.[5]interface {}   �.type..hash.[3]string·f              (type..hash.[3]string   �*type..eq.[3]string·f              $type..eq.[3]string   �:type..hash.[1]interface {}·f              4type..hash.[1]interface {}   �6type..eq.[1]interface {}·f              0type..eq.[1]interface {}   �:type..hash.[2]interface {}·f              4type..hash.[2]interface {}   �6type..eq.[2]interface {}·f              0type..eq.[2]interface {}   ��type..hash.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }·f              �type..hash.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   ��type..eq.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }·f              �type..eq.struct { F uintptr; ctxt *"".Context; p *"".Package; pkga *string; pkgtargetroot string }   ��type..hash.struct { F uintptr; badGoError *error; p *"".Package; name string }·f              �type..hash.struct { F uintptr; badGoError *error; p *"".Package; name string }   ��type..eq.struct { F uintptr; badGoError *error; p *"".Package; name string }·f              �type..eq.struct { F uintptr; badGoError *error; p *"".Package; name string }   �Rtype..hash.struct { a string; b bool }·f              Ltype..hash.struct { a string; b bool }   �Ntype..eq.struct { a string; b bool }·f              Htype..eq.struct { a string; b bool }   �Ztype..hash.[24]struct { a string; b bool }·f              Ttype..hash.[24]struct { a string; b bool }   �Vtype..eq.[24]struct { a string; b bool }·f              Ptype..eq.[24]struct { a string; b bool }   ��go13ld                                                                                                       usr/local/go/pkg/linux_amd64/go/constant.a                                                          0100644 0000000 0000000 00001040516 13101127333 017071  0                                                                                                    ustar 00                                                                0000000 0000000                                                                                                                                                                        !<arch>
__.PKGDEF       0           0     0     644     4504      `
go object linux amd64 go1.6.4 X:none
build id "4cb3e361d5c778548b03e1dd06b866a3ed56b787"

$$
package constant
	import fmt "fmt"
	import math "math"
	import strconv "strconv"
	import utf8 "unicode/utf8"
	import token "go/token"
	import big "math/big"
	type @"".Kind int
	const @"".Unknown @"".Kind = 0x0
	const @"".Bool @"".Kind = 0x1
	const @"".String @"".Kind = 0x2
	const @"".Int @"".Kind = 0x3
	const @"".Float @"".Kind = 0x4
	const @"".Complex @"".Kind = 0x5
	type @"".Value interface { ExactString() (? string); Kind() (? @"".Kind); String() (? string); @"".implementsValue() }
	func @"".MakeUnknown () (? @"".Value) { return (@"".unknownVal{  }) }
	func @"".MakeBool (@"".b·2 bool) (? @"".Value) { return @"".boolVal(@"".b·2) }
	func @"".MakeString (@"".s·2 string "esc:0x12") (? @"".Value) { return @"".stringVal(@"".s·2) }
	func @"".MakeInt64 (@"".x·2 int64) (? @"".Value) { return @"".int64Val(@"".x·2) }
	func @"".MakeUint64 (@"".x·2 uint64) (? @"".Value)
	func @"".MakeFloat64 (@"".x·2 float64) (? @"".Value)
	type @"go/token".Token int
	func (@"go/token".tok·2 @"go/token".Token) IsKeyword () (? bool) { return @"go/token".Token(0x3c) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0x56) }
	func (@"go/token".tok·2 @"go/token".Token) IsLiteral () (? bool) { return @"go/token".Token(0x3) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0xa) }
	func (@"go/token".tok·2 @"go/token".Token) IsOperator () (? bool) { return @"go/token".Token(0xb) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0x3b) }
	func (@"go/token".op·2 @"go/token".Token) Precedence () (? int)
	func (@"go/token".tok·2 @"go/token".Token) String () (? string)
	func @"".MakeFromLiteral (@"".lit·2 string, @"".tok·3 @"go/token".Token, @"".zero·4 uint) (? @"".Value)
	func @"".BoolVal (@"".x·2 @"".Value) (? bool)
	func @"".StringVal (@"".x·2 @"".Value) (? string)
	func @"".Int64Val (@"".x·3 @"".Value) (? int64, ? bool)
	func @"".Uint64Val (@"".x·3 @"".Value) (? uint64, ? bool)
	func @"".Float32Val (@"".x·3 @"".Value) (? float32, ? bool)
	func @"".Float64Val (@"".x·3 @"".Value) (? float64, ? bool)
	func @"".BitLen (@"".x·2 @"".Value) (? int)
	func @"".Sign (@"".x·2 @"".Value) (? int)
	func @"".Bytes (@"".x·2 @"".Value) (? []byte)
	func @"".MakeFromBytes (@"".bytes·2 []byte "esc:0x1") (? @"".Value)
	func @"".Num (@"".x·2 @"".Value) (? @"".Value)
	func @"".Denom (@"".x·2 @"".Value) (? @"".Value)
	func @"".MakeImag (@"".x·2 @"".Value) (? @"".Value)
	func @"".Real (@"".x·2 @"".Value) (? @"".Value)
	func @"".Imag (@"".x·2 @"".Value) (? @"".Value)
	func @"".ToInt (@"".x·2 @"".Value) (? @"".Value)
	func @"".ToFloat (@"".x·2 @"".Value) (? @"".Value)
	func @"".ToComplex (@"".x·2 @"".Value "esc:0x1a") (? @"".Value)
	func @"".UnaryOp (@"".op·2 @"go/token".Token, @"".y·3 @"".Value, @"".prec·4 uint) (? @"".Value)
	func @"".BinaryOp (@"".x·2 @"".Value, @"".op·3 @"go/token".Token, @"".y·4 @"".Value) (? @"".Value)
	func @"".Shift (@"".x·2 @"".Value, @"".op·3 @"go/token".Token, @"".s·4 uint) (? @"".Value)
	func @"".Compare (@"".x·2 @"".Value, @"".op·3 @"go/token".Token, @"".y·4 @"".Value) (? bool)
	func @"".init ()
	type @"".unknownVal struct {}
	func (@"".x·2 @"".unknownVal) ExactString () (? string) { return @"".x·2.String() }
	func (? @"".unknownVal) Kind () (? @"".Kind) { return @"".Kind(0x0) }
	func (? @"".unknownVal) String () (? string) { return string("unknown") }
	func (? @"".unknownVal) @"".implementsValue () {  }
	type @"".boolVal bool
	func (@"".x·2 @"".boolVal) ExactString () (? string) { return @"".x·2.String() }
	func (? @"".boolVal) Kind () (? @"".Kind) { return @"".Kind(0x1) }
	func (@"".x·2 @"".boolVal) String () (? string) { return @"strconv".FormatBool(bool(@"".x·2)) }
	func (? @"".boolVal) @"".implementsValue () {  }
	type @"".stringVal string
	func (@"".x·2 @"".stringVal "esc:0x1") ExactString () (? string)
	func (? @"".stringVal) Kind () (? @"".Kind) { return @"".Kind(0x2) }
	func (@"".x·2 @"".stringVal "esc:0x1") String () (? string)
	func (? @"".stringVal) @"".implementsValue () {  }
	type @"".int64Val int64
	func (@"".x·2 @"".int64Val) ExactString () (? string)
	func (? @"".int64Val) Kind () (? @"".Kind) { return @"".Kind(0x3) }
	func (@"".x·2 @"".int64Val) String () (? string)
	func (? @"".int64Val) @"".implementsValue () {  }
	func @"strconv".FormatBool (@"strconv".b·2 bool) (? string) { if @"strconv".b·2 { return string("true") }; return string("false") }

$$
_go_.o          0           0     0     644     274230    `
go object linux amd64 go1.6.4 X:none

!
  go13ld
fmt.ago/token.amath.amath/big.astrconv.aunicode/utf8.a �$"".unknownVal.Kind      H�D$    �������    "".~r0  type."".Kind   �  Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".boolVal.Kind      H�D$   �������     "".~r0 type."".Kind   �  Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�""".stringVal.Kind      H�D$   ������� 0   "".~r0  type."".Kind   �  Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go� "".int64Val.Kind      H�D$   �������     "".~r0 type."".Kind   �  Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".intVal.Kind      H�D$   �������     "".~r0 type."".Kind   �  Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".ratVal.Kind      H�D$   �������     "".~r0 type."".Kind   �  Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go� "".floatVal.Kind      H�D$   �������     "".~r0 type."".Kind   �  Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�$"".complexVal.Kind      H�D$(   ������� P   "".~r0 @type."".Kind   �  Tgclocals·d0110d631ecd4af0947009e36d46dc99 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�("".unknownVal.String  @  @1�H�    H�\$H�D$   ���������
  &go.string."unknown"       "".~r0  type.string     �   Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�""".boolVal.String  �  �1��D$1�< tH�    H��   H�L$H�D$�H�    H��   ������������    go.string."true"   R  "go.string."false"   0   "".~r0 type.string "".x  type."".boolVal @ @ �@  Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�&"".stringVal.String  �  �dH�%    H;a�E  H��h1�H��$�   H��$�   H�\$pH�$H�\$xH�\$�    H�L$H�D$H�L$HH�$H�D$PH�D$�    H�t$HH�T$PH�\$H��H��   1�1�H�D$8H��E}cH�L$@H��H9���   H)�I��H�� tM�L�D$XL�$H�l$`H�l$�    H�t$HH�T$PH�D$H�L$@H�H�D$8H��H�D$8H��E|�H9�wUH�$    H�t$XH�t$H�L$`H�L$H�    H�\$H�D$    �    H�t$(H�T$0H��$�   H��$�   H��h��    �    ���    ������������������
      z  strconv.Quote   �  <unicode/utf8.RuneCountInString   �  >unicode/utf8.DecodeRuneInString   �  go.string."..."   �  *runtime.concatstring2   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0005  type.string "".autotmp_0003  type.int "".autotmp_0002 type.string "".n _type.int "".i Otype.int "".s ?type.string "".~r0  type.string "".x  "type."".stringVal  ����� � <�)"1HE
  <"�L Tgclocals·f47057354ec566066f8688a4970cff5a Tgclocals·83ead081cd909acab0dcd88a450c1878   @$GOROOT/src/go/constant/value.go�$"".int64Val.String  �  �dH�%    H;av@H�� 1�H�\$0H�\$8H�\$(H�$H�D$
   �    H�L$H�D$H�L$0H�D$8H�� ��    �����������
      d  "strconv.FormatInt   �  0runtime.morestack_noctxt   0@  "".~r0 type.string "".x   type."".int64Val @;? ` �` 
 1/ Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go� "".intVal.String  �  �dH�%    H;av7H��1�H�\$(H�\$0H�\$ H�$�    H�L$H�D$H�L$(H�D$0H����    ����
      R  ,math/big.(*Int).String   �  0runtime.morestack_noctxt   00  "".~r0 type.string "".x  type."".intVal 02/ P �P 
 (( Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go� "".ratVal.String  �  �dH�%    H;avJH�� 1�H�\$0H�\$8H�\$(H�$�    H�D$H�D$H�$�    H�L$H�D$H�L$0H�D$8H�� ��    �
      R  "".rtof   x  $"".floatVal.String   �  0runtime.morestack_noctxt   0@  "".autotmp_0008  type."".floatVal "".~r0 type.string "".x  type."".ratVal @E? ` �` 
 (8 Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·5184031d3a32a42d85027f073f873668   @$GOROOT/src/go/constant/value.go�$"".floatVal.String  �  �dH�%    H�D$�H;A�  H���   1�H��$   H��$  H��$�   �X������ t+H�$�    H�L$H�D$H��$   H��$  H���   �H�D$hH�$�    �D$�D$8H�\$hH�$�    �D$8H�\$H�� ��f(�W�f.�A��@��L!�@8��]  f(�1�H�� |f(��    f.��1  H�� �   f(��    f.���< �  �\$`1�H��$�   H��$�   H��$�   H�� ��   HǄ$�      HǄ$�      H��$�   H�    H�$H�\$`H�\$H�D$    �    H�L$H�D$ H��$�   H�L$pH�H�D$x�=     ufH�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�L$(H�D$0H��$   H��$  H���   �L�CL�$H�D$�    늉����H��$�   W�CCH�\$hH�$H��$�   H�\$�    H�\$H�\$@H��$�   H�$�    �\$H�D$@�H*�f(��    �Y��H,��\$X�    �$H�D$H�H*�f(�f(��\��L$�    H�D$H�T$�\$X�Y�f(�W�W�f.��  W�f.���  ��  W�f(�f(��    f.���  �    f.���  �T$`H�D$P1�H��$�   H��$�   H��$�   H��$�   H��$�   H�� �S  HǄ$�      HǄ$�      H��$�   H�    H�$H�\$`H�\$H�D$    �    H�L$H�D$ H��$�   H�L$pH�H�D$x�=     ��   H�CH�    H�$H�\$PH�\$H�D$    �    H�L$H�D$ H��$�   H��H�L$pH�H�D$x�=     ufH�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�L$(H�D$0H��$   H��$  H���   �L�CL�$H�D$�    �L�CL�$H�D$�    � ���������    �^�H���S����    �Y�f(�H���;���f(������    �Y������1������H��   ������    ����������������B
      �  0math/big.(*Float).String   �  2math/big.(*Float).Float64   �  ,math/big.(*Float).Sign   �  *$f64.7fefffffffffffff   �  *$f64.ffefffffffffffff   �  type.float64   �  runtime.convT2E   � (runtime.writeBarrier   �   go.string."%.6g"   �  fmt.Sprintf   �  .runtime.writebarrierptr   �	  2math/big.(*Float).MantExp   �	  2math/big.(*Float).Float64   �
  *$f64.3fd34413509f79ff   �
  *$f64.4024000000000000   �  math.Pow   �  *$f64.3feffffef39085f5   �  *$f64.4024000000000000   �  type.float64   �  runtime.convT2E   � (runtime.writeBarrier   �  type.int64   �  runtime.convT2E   � (runtime.writeBarrier   �  (go.string."%.6ge%+d"   �  fmt.Sprintf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  *$f64.4024000000000000   �  *$f64.4024000000000000   �  *$f64.bff0000000000000   �  0runtime.morestack_noctxt   0�  2"".autotmp_0036  "type.interface {} "".autotmp_0035  "type.interface {} "".autotmp_0034 �(type.[2]interface {} "".autotmp_0031  &type.[]interface {} "".autotmp_0030  type.float64 "".autotmp_0029 �"type.interface {} "".autotmp_0028 �(type.[1]interface {} "".autotmp_0025 �&type.[]interface {} "".autotmp_0024  type.bool "".autotmp_0022  type.string "".autotmp_0021 �type.int64 "".autotmp_0020  type.float64 "".autotmp_0019  type.int64 "".autotmp_0018  type.float64 "".autotmp_0016  type.float64 "".autotmp_0014 �type.float64 "".autotmp_0013  type.string "".autotmp_0012 �type.float64 "".e �type.int64 "".exp �type.int "".mant O&type.math/big.Float "".x �type.float64 "".f �(type.*math/big.Float "".~r0 type.string "".x   type."".floatVal <�S���������� �
 n�1+
��%M*
�) 2 L0�l4:��4� Tgclocals·948c285cf1025b717e2658a3cccfd415 Tgclocals·ec147618165580e6a5d760bf3329b6ac   @$GOROOT/src/go/constant/value.go�("".complexVal.String  �  �dH�%    H;a�t  H��   1�H��$�   H��$�   1�H�\$`H�\$hH�\$pH�\$xH�\$`H�� �/  H�D$P   H�D$X   H�\$HH��$�   H�H�$H�KH�L$�    H�L$H�D$H�\$HH�L$8H�H�D$@�=     ��   H�CH��$�   H�H�$H�KH�L$�    H�L$H�D$H�\$HH��H�L$8H�H�D$@�=     u]H�CH�    H�$H�D$
   H�\$HH�\$H�\$PH�\$H�\$XH�\$ �    H�L$(H�D$0H��$�   H��$�   H�Ā   �L�CL�$H�D$�    �L�CL�$H�D$�    �2����������    �o������������������
      �  runtime.convI2E   � (runtime.writeBarrier   �  runtime.convI2E   � (runtime.writeBarrier   �  ,go.string."(%s + %si)"   �  fmt.Sprintf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   `�  "".autotmp_0043  "type.interface {} "".autotmp_0042 �"type.interface {} "".autotmp_0041 ?(type.[2]interface {} "".autotmp_0038 o&type.[]interface {} "".~r0 @type.string "".x  $type."".complexVal  ����2� � 
��  ��4> Tgclocals·23322ef3fd8702babe318da8c8d339e7 Tgclocals·341b909b97472a89efab32cbd0761e34   @$GOROOT/src/go/constant/value.go�2"".unknownVal.ExactString  @  @1�1�H�    H��   H�\$H�D$����  &go.string."unknown"       "".~r0  type.string "".x  $type."".unknownVal     �   Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�,"".boolVal.ExactString  �  �1��D$1�1�< tH�    H��   H�L$H�D$�H�    H��   ����������$   go.string."true"   V  "go.string."false"   0   "".~r0 type.string "".x  type."".boolVal @ @ �@  Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�0"".stringVal.ExactString  �  �dH�%    H;avAH�� 1�H�\$8H�\$@H�\$(H�$H�\$0H�\$�    H�L$H�D$H�L$8H�D$@H�� ��    ����������
      f  strconv.Quote   �  0runtime.morestack_noctxt   @@  "".~r0  type.string "".x  "type."".stringVal @<? ` �` 
 2. Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�."".int64Val.ExactString  �  �dH�%    H;av7H��1�H�\$(H�\$0H�\$ H�$�    H�L$H�D$H�L$(H�D$0H����    ����
      R  $"".int64Val.String   �  0runtime.morestack_noctxt   00  "".~r0 type.string "".x   type."".int64Val 02/ P �P 
 (( Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�*"".intVal.ExactString  �  �dH�%    H;av7H��1�H�\$(H�\$0H�\$ H�$�    H�L$H�D$H�L$(H�D$0H����    ����
      R   "".intVal.String   �  0runtime.morestack_noctxt   00  "".~r0 type.string "".x  type."".intVal 02/ P �P 
 (( Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�*"".ratVal.ExactString  �  �dH�%    H;a��   H�� 1�H�\$0H�\$8H�D$(H�D$H�$�    H�L$�\$�� t,H�� t"H�$�    H�L$H�D$H�L$0H�D$8H�� É��H�$�    H�L$H�D$H�L$0H�D$8H�� ��    �c������

      d  *math/big.(*Rat).IsInt   �  ,math/big.(*Int).String   �  ,math/big.(*Rat).String   �  0runtime.morestack_noctxt   0@  "".autotmp_0051  type.string "".r $type.*math/big.Rat "".~r0 type.string "".x  type."".ratVal @U?@%? � �#,"	  1Q Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·0c8aa8e80191a30eac23f1a218103f16   @$GOROOT/src/go/constant/value.go�."".floatVal.ExactString  �  �dH�%    H;avEH��(1�H�\$8H�\$@H�\$0H�$�D$pH�D$    �    H�L$H�D$ H�L$8H�D$@H��(��    ������
      n  ,math/big.(*Float).Text   �  0runtime.morestack_noctxt   0P  "".~r0 type.string "".x   type."".floatVal P@O ` �` 
 6* Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�2"".complexVal.ExactString  �  �dH�%    H�D$�H;A�  H��   1�H��$�   H��$�   H��$�   H��$�   H�D$@H�$H�L$8H�Y ��H�\$H�\$hH�\$H�\$pH��$�   H��$�   H�D$@H�$H�L$8H�Y ��H�\$H�\$XH�\$H�\$`1�H��$�   H��$�   H��$�   H��$�   H��$�   H�� �G  HǄ$�      HǄ$�      H�\$xH�    H�$H�\$hH�\$H�D$    �    H�L$H�D$ H�\$xH�L$HH�H�D$P�=     ��   H�CH�    H�$H�\$XH�\$H�D$    �    H�L$H�D$ H�\$xH��H�L$HH�H�D$P�=     ucH�CH�    H�$H�D$
   H�\$xH�\$H��$�   H�\$H��$�   H�\$ �    H�L$(H�D$0H��$�   H��$�   H�İ   �L�CL�$H�D$�    �L�CL�$H�D$�    �&���������    ��������
      �       �       �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  type.string   �  runtime.convT2E   � (runtime.writeBarrier   �  ,go.string."(%s + %si)"   �  fmt.Sprintf   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   `�  "".autotmp_0062  "type.interface {} "".autotmp_0061 �"type.interface {} "".autotmp_0060 ?(type.[2]interface {} "".autotmp_0057 o&type.[]interface {} "".autotmp_0055 �type.string "".autotmp_0054 �type.string "".~r0 @type.string "".x  $type."".complexVal  ����2� � �1�  S8��42 Tgclocals·ae0b17ff166fa616635ce4bad0c70f06 Tgclocals·a19b4fb8a607611184c7491e4d9543cb   @$GOROOT/src/go/constant/value.go�:"".unknownVal.implementsValue      ����������������        �  Tgclocals·33cdeccccebe80329f1fdbee7f5874cb Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�4"".boolVal.implementsValue      ����������������       �  Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�8"".stringVal.implementsValue      ����������������        �  Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�6"".int64Val.implementsValue      ����������������       �  Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�2"".ratVal.implementsValue      ����������������       �  Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�2"".intVal.implementsValue      ����������������       �  Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�6"".floatVal.implementsValue      ����������������       �  Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�:"".complexVal.implementsValue      ���������������� @      �  Tgclocals·31b2ddfd7c7062d584469c95698a3e1d Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".newInt  �  �dH�%    H;av#H��H�    H�$�    H�\$H�\$H����    ���������
      ,  "type.math/big.Int   >  "runtime.newobject   f  0runtime.morestack_noctxt      "".~r0  $type.*math/big.Int   @ �@ 
 " Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".newRat  �  �dH�%    H;av#H��H�    H�$�    H�\$H�\$H����    ���������
      ,  "type.math/big.Rat   >  "runtime.newobject   f  0runtime.morestack_noctxt      "".~r0  $type.*math/big.Rat   @ �@ 
 " Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".newFloat  �  �dH�%    H;av:H��H�    H�$�    H�\$H�$H�D$   �    H�\$H�\$ H����    �

      ,  &type.math/big.Float   >  "runtime.newobject   l  2math/big.(*Float).SetPrec   �  0runtime.morestack_noctxt   0  "".autotmp_0068  (type.*math/big.Float "".~r0  (type.*math/big.Float 05/ P �P 
 2 Tgclocals·5184031d3a32a42d85027f073f873668 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".i64toi  �  �dH�%    H;avDH��1�H�\$(H�    H�$�    H�\$H�$H�\$ H�\$�    H�D$1�H�D$(H����    �������

      :  "type.math/big.Int   L  "runtime.newobject   |  0math/big.(*Int).SetInt64   �  0runtime.morestack_noctxt    0  "".autotmp_0070  $type.*math/big.Int "".~r1 type."".intVal "".x   type."".int64Val 0?/ ` �` 
 %; Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".i64tor  �  �dH�%    H;avDH��1�H�\$(H�    H�$�    H�\$H�$H�\$ H�\$�    H�D$1�H�D$(H����    �������

      :  "type.math/big.Rat   L  "runtime.newobject   |  0math/big.(*Rat).SetInt64   �  0runtime.morestack_noctxt    0  "".autotmp_0073  $type.*math/big.Rat "".~r1 type."".ratVal "".x   type."".int64Val 0?/ ` �` 
 %; Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".i64tof  �  �dH�%    H;av8H��1�H�\$(�    H�$H�$H�\$ H�\$�    H�D$1�H�D$(H����    ���
      6  "".newFloat   d  4math/big.(*Float).SetInt64   �  0runtime.morestack_noctxt    0  "".autotmp_0076  (type.*math/big.Float "".~r1  type."".floatVal "".x   type."".int64Val 03/
 P �P 
 6 Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".itor  �  �dH�%    H;avDH��1�H�\$(H�    H�$�    H�\$H�$H�\$ H�\$�    H�D$1�H�D$(H����    �������

      :  "type.math/big.Rat   L  "runtime.newobject   |  ,math/big.(*Rat).SetInt   �  0runtime.morestack_noctxt    0  "".autotmp_0079  $type.*math/big.Rat "".~r1 type."".ratVal "".x  type."".intVal 0?/ ` �` 
 %; Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".itof  �  �dH�%    H;av8H��1�H�\$(�    H�$H�$H�\$ H�\$�    H�D$1�H�D$(H����    ���
      6  "".newFloat   d  0math/big.(*Float).SetInt   �  0runtime.morestack_noctxt    0  "".autotmp_0082  (type.*math/big.Float "".~r1  type."".floatVal "".x  type."".intVal 03/
 P �P 
 6 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".rtof  �  �dH�%    H;a��   H��01�H�\$@�    H�$H�D$8H�� tzH�$H�D$�    H�\$H�\$(�    H�$H�\$ H�\$8H�$�    H�D$H�\$ H�$H�D$�    H�L$(H�D$H�$H�L$H�D$�    H�D$1�H�D$@H��0É ��    �F���������
      >  "".newFloat   x  0math/big.(*Float).SetInt   �  "".newFloat   �  *math/big.(*Rat).Denom   �  0math/big.(*Float).SetInt   �  *math/big.(*Float).Quo   �  0runtime.morestack_noctxt    `  "".autotmp_0087  (type.*math/big.Float "".autotmp_0086  $type.*math/big.Int "".autotmp_0085  (type.*math/big.Float "".autotmp_0084 (type.*math/big.Float "".a (type.*math/big.Float "".~r1  type."".floatVal "".x  type."".ratVal `�_`_ � �,>$  ,* Tgclocals·f7309186bf9eeb0f8ece2eb16f2dc110 Tgclocals·b40f0f67eae216e69d0bb41a8427b144   @$GOROOT/src/go/constant/value.go�"".vtoc  �  �dH�%    H;a��   H��`1�H�\$xH��$�   H��$�   H��$�   H�D$8    1�H�\$@H�\$HH�\$PH�\$XH�\$hH�\$@H�\$pH�\$HH�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�l$PH�H�M H�KH�MH�\$@H�\$xH�\$HH��$�   H�\$PH��$�   H�\$XH��$�   H��`��    �������
      �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   `�  "".autotmp_0091 ?$type."".complexVal "".autotmp_0090 O type."".int64Val "".~r1  $type."".complexVal "".x  type."".Value ��� � 
��  �a Tgclocals·aa5118865dd28fc3eaacbfc830efb456 Tgclocals·4cf9735ef08c57d91ff7cf30faacc15b   @$GOROOT/src/go/constant/value.go�"".makeInt  �  �dH�%    H;a�i  H��`1�H�\$pH�\$xH�    H�$H�\$hH�\$�    H�L$hH�\$H�� ��   H�$H�    H�\$�    H�L$hH�\$H�� ��   H�� ��   H�qH�t$HH�QH�iH�l$XH�T$PH�� uf1���� tH��H�D$8H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$pH�\$0H�\$xH��`�H�� vH���    ��`���1�H�L$@H�    1�H9�tH�\$@H�\$xH�D$pH��`�H�    H�$H�    H�\$H�    H�\$�    H�D$��    �z������������� 
      L  "".minInt64   r  &math/big.(*Int).Cmp   �  "".maxInt64   �  &math/big.(*Int).Cmp   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $runtime.panicindex   �  4go.itab."".intVal."".Value   �  type."".intVal   �  type."".Value   �  4go.itab."".intVal."".Value   �   runtime.typ2Itab   �  0runtime.morestack_noctxt   0�  "".autotmp_0098 ?type."".intVal "".autotmp_0097 O type."".int64Val "".autotmp_0095  type.int math/big.z·2 /"type.math/big.nat "".~r1 type."".Value "".x  $type.*math/big.Int ,����A��/� � �#W�X  8�  Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·83ead081cd909acab0dcd88a450c1878   @$GOROOT/src/go/constant/value.go�"".makeRat  �  �dH�%    H;a��  H��HH�L$P1�H�\$XH�\$`H�� �i  H�L$@H�$�    H�\$H�\$(H�\$@H�$�    H�\$H��   }yH�\$(H�$�    H�\$H��   }]1�H�\$PH�\$8H�    1�H9�tH�\$8H�\$`H�D$XH��H�H�    H�$H�    H�\$H�    H�\$�    H�D$��    H�$H�$H�\$@H�\$�    H�\$H�\$ �    H�$H�$H�\$(H�\$�    H�L$ H�D$H�$H�L$H�D$�    H�D$1�H�D$0H�    1�H9�tH�\$0H�\$`H�D$XH��H�H�    H�$H�    H�\$H�    H�\$�    H�D$뽉�����    �T�������(
      x  *math/big.(*Rat).Denom   �  ,math/big.(*Int).BitLen   �  ,math/big.(*Int).BitLen   �  4go.itab."".ratVal."".Value   �  type."".ratVal   �  type."".Value   �  4go.itab."".ratVal."".Value   �   runtime.typ2Itab   �  "".newFloat   �  0math/big.(*Float).SetInt   �  "".newFloat   �  0math/big.(*Float).SetInt   �  *math/big.(*Float).Quo   �  8go.itab."".floatVal."".Value   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  0runtime.morestack_noctxt   0�  "".autotmp_0110  type.*uint8 "".autotmp_0107 / type."".floatVal "".autotmp_0106  (type.*math/big.Float "".autotmp_0105  (type.*math/big.Float "".autotmp_0103 type."".ratVal 
"".fa O(type.*math/big.Float "".b ?$type.*math/big.Int "".a $type.*math/big.Int "".~r1 type."".Value "".x  $type.*math/big.Rat .�������6� � ,�(8]&&p , ;�V! Tgclocals·add78ec634cef78099972ccd9d767bc6 Tgclocals·549df0c0b9c1ff589e7323390661782b   @$GOROOT/src/go/constant/value.go�"".makeFloat  �  �dH�%    H;a��   H��(1�H�\$8H�\$@H�\$0H�$�    H�\$H�� uSH�    1�H9�tH�    H�\$@H�D$8H��(�H�    H�$H�    H�\$H�    H�\$�    H�D$�1�H�\$0H�\$ H�    1�H9�tH�\$ H�\$@H�D$8H��(�H�    H�$H�    H�\$H�    H�\$�    H�D$��    �
�������������
      Z  ,math/big.(*Float).Sign   ~  8go.itab."".floatVal."".Value   �  "".floatVal0   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  8go.itab."".floatVal."".Value   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  0runtime.morestack_noctxt   0P  "".autotmp_0116  type.*uint8 "".autotmp_0114  type."".floatVal "".~r1 type."".Value "".x  (type.*math/big.Float PHOP\OP/O � �#S]	  ,�  Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·0c8aa8e80191a30eac23f1a218103f16   @$GOROOT/src/go/constant/value.go�"".makeComplex  �  �dH�%    H;a��   H��X1�H��$�   H��$�   1�H�\$8H�\$@H�\$HH�\$PH�\$`H�\$8H�\$hH�\$@H�\$pH�\$HH�\$xH�\$PH�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H��$�   H�\$0H��$�   H��X��    �5��������
      �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   `�  "".autotmp_0119 ?$type."".complexVal "".~r2 @type."".Value 
"".im  type."".Value 
"".re  type."".Value ��� � �)�  �3 Tgclocals·8c2f8f990ab0a90930a640c5478081b4 Tgclocals·4cf9735ef08c57d91ff7cf30faacc15b   @$GOROOT/src/go/constant/value.go�."".makeFloatFromLiteral  �  �dH�%    H;a�,  H��81�H�\$PH�\$X�    H�$H�$H�\$@H�\$H�\$HH�\$�    H�L$�\$ �� ��   H�L$(H�$�    �\$�� ��   H�    H�$�    H�\$H�$H�\$@H�\$H�\$HH�\$�    H�D$1�H�D$0H�    1�H9�tH�\$0H�\$XH�D$PH��8�H�    H�$H�    H�\$H�    H�\$�    H�D$�H�\$(H�$�    H�L$H�D$H�L$PH�D$XH��8�1�H�\$PH�\$XH��8��    �����������
      H  "".newFloat   �  6math/big.(*Float).SetString   �  "".smallRat   �  "type.math/big.Rat   �  "runtime.newobject   �  2math/big.(*Rat).SetString   �  4go.itab."".ratVal."".Value   �  type."".ratVal   �  type."".Value   �  4go.itab."".ratVal."".Value   �   runtime.typ2Itab   �  "".makeFloat   �  0runtime.morestack_noctxt   @p  "".autotmp_0123 type."".ratVal "".f (type.*math/big.Float "".~r1  type."".Value "".lit  type.string  p�opUopo � $�#97X'  #Bx@ Tgclocals·55cc6ee7528f0b48e5a6d9bfba36524a Tgclocals·e48b749e068cae7c3a399141c10fe5f0   @$GOROOT/src/go/constant/value.go�"".smallRat  �  �dH�%    H;avWH��H�L$ �Y����< u6H�$H�D$    �    H�D$H= ���~H=   �D$(H����D$( ���D$( H����    ����
      h  2math/big.(*Float).MantExp   �  0runtime.morestack_noctxt    0  "".~r1 type.bool "".x  (type.*math/big.Float 0A/0/ p �
	
 
 3= Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".MakeUnknown  �  �dH�%    H;avfH��81�H�\$@H�\$H1�H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$@H�\$0H�\$HH��8��    �����
      H  $type."".unknownVal   ^  type."".Value   v  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt    p  "".autotmp_0128  $type."".unknownVal "".~r0  type."".Value pao � 
�� 
 W) Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".MakeBool  �  �dH�%    H;avmH��@1�H�\$PH�\$X�\$H�\$?H�    H�$H�    H�\$H�    H�\$H�\$?H�\$H�D$     �    H�\$(H�\$PH�\$0H�\$XH��@��    �z�������������
      V  type."".boolVal   l  type."".Value   �  6go.itab."".boolVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   0�  "".autotmp_0129 type."".boolVal "".~r1 type."".Value "".b  type.bool �h � 
�� 
 ^2 Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".MakeString  �  �dH�%    H;avxH��H1�H�\$`H�\$hH�\$PH�\$8H�\$XH�\$@H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$`H�\$0H�\$hH��H��    �o������������������
      l  "type."".stringVal   �  type."".Value   �  :go.itab."".stringVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   @�  "".autotmp_0130 "type."".stringVal "".~r1  type."".Value "".s  type.string �s� � 
�� 
 i7 Tgclocals·f47057354ec566066f8688a4970cff5a Tgclocals·d8fdd2a55187867c76648dc792366181   @$GOROOT/src/go/constant/value.go�"".MakeInt64  �  �dH�%    H;avnH��@1�H�\$PH�\$XH�\$HH�\$8H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$PH�\$0H�\$XH��@��    �y������������
      X   type."".int64Val   n  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   0�  "".autotmp_0131  type."".int64Val "".~r1 type."".Value "".x  type.int64 �i � 
�� 
 _1 Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".MakeUint64  �  �dH�%    H;a�  H��HH�D$P1�H�\$XH�\$`H�       �H9�sYH�D$8H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$XH�\$0H�\$`H��H�H�    H�$�    H�\$H�$H�\$PH�\$�    H�D$1�H�D$@H�    1�H9�tH�\$@H�\$`H�D$XH��H�H�    H�$H�    H�\$H�    H�\$�    H�D$��    ������
      ~   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "type.math/big.Int   �  "runtime.newobject   �  2math/big.(*Int).SetUint64   �  4go.itab."".intVal."".Value   �  type."".intVal   �  type."".Value   �  4go.itab."".intVal."".Value   �   runtime.typ2Itab   �  0runtime.morestack_noctxt   0�  
"".autotmp_0135 type."".intVal "".autotmp_0134  $type.*math/big.Int "".autotmp_0132  type."".int64Val "".~r1 type."".Value "".x  type.uint64 *�x��U��/� � �(Y�  r� Tgclocals·f56b2291fa344104975cb6587be42b9b Tgclocals·0c8aa8e80191a30eac23f1a218103f16   @$GOROOT/src/go/constant/value.go�"".MakeFloat64  �  �dH�%    H;a��  H��H�\$P1�H�\$XH�\$`f(�1�H�� |�    f.���  H�� �q  �    f.���< �  f.�����H	�< ��   W�f.�u_z]H�D$8    H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$XH�\$0H�\$`H��H�H�    H�$�    H�\$H�$�D$P�D$�    H�D$1�H�D$@H�    1�H9�tH�\$@H�\$`H�D$XH��H�H�    H�$H�    H�\$H�    H�\$�    H�D$�1�H�    H�$H�    H�\$H�    H�\$H�\$8H�\$H�D$     �    H�\$(H�\$XH�\$0H�\$`H��H�1�����H��   �����    �!����(
      r  *$f64.7fefffffffffffff   �  *$f64.ffefffffffffffff   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "type.math/big.Rat   �  "runtime.newobject   �  4math/big.(*Rat).SetFloat64   �  4go.itab."".ratVal."".Value   �  type."".ratVal   �  type."".Value   �  4go.itab."".ratVal."".Value   �   runtime.typ2Itab   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   0�  "".autotmp_0144  type.bool "".autotmp_0142 type."".ratVal "".autotmp_0141  $type.*math/big.Rat "".autotmp_0139  type."".int64Val "".autotmp_0138 $type."".unknownVal "".~r1 type."".Value "".x  type.float64 :����W������ � &�)T]�V  ��D< Tgclocals·f56b2291fa344104975cb6587be42b9b Tgclocals·0c8aa8e80191a30eac23f1a218103f16   @$GOROOT/src/go/constant/value.go�$"".MakeFromLiteral  �  �dH�%    H��$����H;A��  H��  H��$�  H��$�  H��$�  1�H��$�  H��$�  H��$�  H�� t]H�    H��$h  HǄ$p  2   H�    H�$H��$h  H�\$H�D$    �    H�\$H�H�$H�KH�L$�    H���m  H����  H�$H�D$H�D$    H�D$@   �    H�D$ H�L$(H�\$0H��$   H��$�   H�� ubH�D$HH�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�İ  �H�    H�$�    H�\$H�$H��$�  H�\$H��$�  H�\$H�D$    �    H�L$ �\$(�� ta1�H�L$PH�    1�H9�tH�\$PH��$�  H��$�  H�İ  �H�    H�$H�    H�\$H�    H�\$�    H�D$�1�H�    H�$H�    H�\$H�    H�\$H�\$@H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�İ  �H��uJH�$H�D$�    H�D$H�L$H��$�   H��$�   H�� �i���H��$�  H��$�  H�İ  �H�l$@1�H��$(  H��$0  H��$(  H�� �,  HǄ$�     HǄ$�     H��$x  H�    H�$H�\$@H�\$H�D$    �    H�L$H�D$ H��$x  H��$  H�H��$   �=     ��   H�CH�    H�$H�D$   H��$x  H�\$H��$�  H�\$H��$�  H�\$ �    H�\$(H��$h  H�\$0H��$p  H�    H�$H��$h  H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M���������H����  H�� �����H��H��H9���  H�*���i�����H��H��H9��~  H��$X  H�$H��$`  H�\$�    H�D$H�\$H��$�   H��$�   H�� �q���H�D$H    H�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�l$(H�T$0H��$8  H��$@  H��$�   H��$�   1�H�\$XH�\$`1�H��$�  H��$�  H��$�  H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$�  H��$�  H�İ  ��    �    H����   H������H��H��H9���   H����   H��H��H�� tH��H��$X  H�,$H��$`  H�\$�D$'�    �D$H�L$0H�\$8H��$�   H��$�   H�� �����Hc�H��1�H�\$hH�\$pH�D$HH�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�L$(H�D$0H��$�  H��$�  H�İ  ��    H��	�����H�$H�D$�    H�L$H��$�   H�T$H��$�   H�D$ H�\$(H��$  H��$  H�� �����1�H�\$xH��$�   H��$�   H��$H  H��$�   H��$P  H�    H�$H�    H�\$H�    H�\$H��$H  H�\$H�D$     �    H�L$(H�D$0H��$�  H��$�  H�İ  ��    �������n
      �  |go.string."MakeFromLiteral called with non-zero last argument"   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �   strconv.ParseInt   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "type.math/big.Int   �  "runtime.newobject   �  2math/big.(*Int).SetString   �  4go.itab."".intVal."".Value   �  type."".intVal   �  type."".Value   �  4go.itab."".intVal."".Value   �   runtime.typ2Itab   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �	  runtime.convT2I   �
  ."".makeFloatFromLiteral   �  &type.go/token.Token   �  runtime.convT2E   � (runtime.writeBarrier   �  Fgo.string."%v is not a valid token"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  ."".makeFloatFromLiteral   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �  $runtime.panicslice   �  $runtime.panicindex   �  &strconv.UnquoteChar   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $runtime.panicslice   �  strconv.Unquote   �  "type."".stringVal   �  type."".Value   �  :go.itab."".stringVal."".Value   �  runtime.convT2I   �  0runtime.morestack_noctxt   `�  H"".autotmp_0173 �"type.interface {} "".autotmp_0172 �(type.[1]interface {} "".autotmp_0169 o&type.[]interface {} "".autotmp_0168  type."".Value "".autotmp_0167  type."".Value "".autotmp_0165  type."".Value "".autotmp_0164 �type."".Value "".autotmp_0161 �$type."".unknownVal "".autotmp_0160  type.string "".autotmp_0159 �&type.go/token.Token "".autotmp_0158 �"type."".stringVal "".autotmp_0157   type."".int64Val "".autotmp_0156  type.string "".autotmp_0155  type.int "".autotmp_0154 ?$type."".complexVal "".autotmp_0153   type."".int64Val "".autotmp_0152 �type.string "".autotmp_0150 �type."".intVal "".autotmp_0148 � type."".int64Val "".autotmp_0147 �type.string "".~r1 �type."".Value "".s �type.string "".~r1 �type."".Value "".~r2 �type."".Value 
"".im �type."".Value 
"".re �type."".Value "".err �type.error "".s �type.string "".err �type.error 
"".im �type."".Value "".x �type."".Value "".err �type.error "".~r3 @type."".Value "".zero 0type.uint "".tok  &type.go/token.Token "".lit  type.string f"����������O���������� � ~�L]

EbPa>_72.�'
)Q�

st

L�E D �P�D�v@.lh�'�
4 Tgclocals·03a89d916197104e2ad001cc20167921 Tgclocals·e6d79eb2ebb897d590c99339e042c95b   @$GOROOT/src/go/constant/value.go�"".BoolVal  �	  �	dH�%    H�D$�H;A�-  H��   H��$�   H��$�   H�L$pH�$H�D$xH�D$�    �L$�L$<����
&uU�D$; H�    H�$H�\$pH�\$H�\$xH�\$H�\$;H�\$�    �L$<�\$ �� t�\$;��$�   H�Ĩ   Á��|~?uJ1�H�    H�$H�\$pH�\$H�\$xH�\$H�\$;H�\$�    �\$ �� tƄ$�    H�Ĩ   �H�T$pH�L$x1�H�\$`H�\$hH�\$`H�� �  HǄ$�      HǄ$�      H��$�   H�T$@H�$H�L$HH�L$�    H�L$H�D$H��$�   H�L$PH�H�D$X�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    �����
      �  $runtime.ifacethash   �  type."".boolVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  2go.string."%v not a Bool"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �	  0runtime.morestack_noctxt   0�  "".autotmp_0183 �"type.interface {} "".autotmp_0182 �(type.[1]interface {} "".autotmp_0179 /&type.[]interface {} "".autotmp_0178 �type.uint32 "".autotmp_0176 otype."".Value "".autotmp_0175 Otype.string "".x �type."".Value "".x �$type."".unknownVal "".x �type."".boolVal "".~r1  type.bool "".x  type."".Value .����Q���� � &�yB
�  B�p@. Tgclocals·aa52d274abdec77c8c6f0039727529fb Tgclocals·60492e1505747e8ca36c9c8f244a1b59   @$GOROOT/src/go/constant/value.go�"".StringVal  �
  �
dH�%    H�D$�H;A�~  H��   W�D$P1�H��$�   H��$�   H��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$�L$<���|~?u^1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� t1�H��$�   H��$�   H�ĸ   Á��n�ul1�H�\$PH�\$XH�    H�$H��$�   H�\$H��$�   H�\$H�\$PH�\$�    �\$ �� t"H�\$PH��$�   H�\$XH��$�   H�ĸ   �H��$�   H��$�   1�H�\$pH�\$xH�\$pH�� �  HǄ$�      HǄ$�      H��$�   H�T$@H�$H�L$HH�L$�    H�L$H�D$H��$�   H�L$`H�H�D$h�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    �`���
      �  $runtime.ifacethash   �  $type."".unknownVal   �  $runtime.assertI2T2   �  "type."".stringVal   �  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  6go.string."%v not a String"   �  fmt.Sprintf   �  type.string   �	  runtime.convT2E   �	  runtime.gopanic   �
  .runtime.writebarrierptr   �
  0runtime.morestack_noctxt   @�  "".autotmp_0192 �"type.interface {} "".autotmp_0191 �(type.[1]interface {} "".autotmp_0188 /&type.[]interface {} "".autotmp_0187 �type.uint32 "".autotmp_0185 otype."".Value "".autotmp_0184 Otype.string "".x �type."".Value "".x �$type."".unknownVal "".x �"type."".stringVal "".~r1  type.string "".x  type."".Value .����s����
 � (�9�R"�
  b�p@. Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc Tgclocals·29c773ae5a332cdcf56287cee2ea280d   @$GOROOT/src/go/constant/value.go�"".Int64Val  �  �dH�%    H�D$�H;A�  H��   1�H�D$HH��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$�L$<���TuhH�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �L$<�\$ �� tH�\$@H��$�   Ƅ$�   H�ĸ   Á��|~?u`1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tHǄ$�       Ƅ$�    H�ĸ   Á�@��q��   1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �\$ �� tXH�L$HH�� tIH�qH�AH�iH�� u%1���� tH��H��$�   Ƅ$�    H�ĸ   �H�� vH����    ��H��$�   H��$�   1�H�\$pH�\$xH�\$pH�� �  HǄ$�      HǄ$�      H��$�   H�T$PH�$H�L$XH�L$�    H�L$H�D$H��$�   H�L$`H�H�D$h�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    �����������������$
      �  $runtime.ifacethash   �   type."".int64Val   �  $runtime.assertI2T2   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  $runtime.panicindex   �  runtime.convI2E   �	 (runtime.writeBarrier   �	  2go.string."%v not an Int"   �
  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   @�  "".autotmp_0204 �"type.interface {} "".autotmp_0203 �(type.[1]interface {} "".autotmp_0200 /&type.[]interface {} "".autotmp_0199 �type.uint32 "".autotmp_0197 otype."".Value "".autotmp_0196 Otype.string "".autotmp_0194  type.int "".x �type."".Value "".x �$type."".unknownVal "".x �type."".intVal "".x � type."".int64Val "".~r2 0type.bool "".~r1  type.int64 "".x  type."".Value <����g������� � 0�&�LQX�   O�ip@.' Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·1170e30e7a2c29fab9e9231402d8c543   @$GOROOT/src/go/constant/value.go�"".Uint64Val  �  �dH�%    H�D$�H;A��  H���   1�H�D$HH��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$�L$<���TuqH�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �L$<�\$ �� t&H�\$@H��$�   H�\$@H�� ��$�   H���   Á��|~?u`1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tHǄ$�       Ƅ$�    H���   Á�@��q�
  1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �\$ �� ��   H�\$HH�� ��   H�SH��$�   H�KH�kH��$�   H��$�   H�� uo1�H��H�D$HH�hH�� uA1�H��$�   H�� |'H�\$HH�$�    H�\$H��@��$�   H���   �Ƅ$�    ����� t	H�������H��   �H�� vH���    ��N���H��$�   H��$�   1�H�\$pH�\$xH�\$pH�� �  HǄ$�      HǄ$�      H��$�   H�T$PH�$H�L$XH�L$�    H�L$H�D$H��$�   H�L$`H�H�D$h�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    �V���������&
      �  $runtime.ifacethash   �   type."".int64Val   �  $runtime.assertI2T2   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  ,math/big.(*Int).BitLen   �	  $runtime.panicindex   �
  runtime.convI2E   � (runtime.writeBarrier   �  2go.string."%v not an Int"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   @�  $"".autotmp_0219 �"type.interface {} "".autotmp_0218 �(type.[1]interface {} "".autotmp_0215 /&type.[]interface {} "".autotmp_0214  type.uint64 "".autotmp_0213 �type.uint32 "".autotmp_0211 �type."".Value "".autotmp_0210 type.string "".autotmp_0209  type.int "".autotmp_0208  type.int "".autotmp_0206  type.int math/big.z·2 _"type.math/big.nat "".x �type."".Value "".x �$type."".unknownVal "".x �type."".intVal "".x � type."".int64Val "".~r2 0type.bool "".~r1  type.uint64 "".x  type."".Value <����g������� � 2�&�&LU�� " O��p@.! Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·50c543803d8632f8d2f7062c2b1cdc18   @$GOROOT/src/go/constant/value.go�"".Float32Val  �  �dH�%    H�D$�H;A�H  H���   W�D$HD$PW�H��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$���T�_  �L$<��1��u~1�H�\$XH�    H�$H��$�   H�\$H��$�   H�\$H�\$XH�\$�    �L$<�\$ �� t5H�\$XH�$�    �D$�\$��$�   �� ��$�   H���   Á��TuwH�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �\$ �� t0H�\$@�H*���$�   H�l$@�H,�H9���$�   H���   �H��$�   H��$�   1�H��$�   H��$�   H��$�   H�� �  HǄ$�      HǄ$�      H��$�   H�T$`H�$H�L$hH�L$�    H�L$H�D$H��$�   H�L$pH�H�D$x�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<����>uz1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �L$<�\$ �� t1H�\$HH�$�    �D$�\$��$�   ��$�   H���   Á��|~?u`1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tW���$�   Ƅ$�    H���   Á�@��q�����1�H�\$PH�    H�$H��$�   H�\$H��$�   H�\$H�\$PH�\$�    �\$ �� �g����    H�$H�$H�\$PH�\$�    H�\$H�$�    �D$�\$��$�   �� ��$�   H���   ��    ����������4
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  2math/big.(*Float).Float32   �   type."".int64Val   �  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  4go.string."%v not a Float"   �	  fmt.Sprintf   �	  type.string   �
  runtime.convT2E   �
  runtime.gopanic   �
  .runtime.writebarrierptr   �  type."".ratVal   �  $runtime.assertI2T2   �  .math/big.(*Rat).Float32   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  "".newFloat   �  0math/big.(*Float).SetInt   �  2math/big.(*Float).Float32   �  0runtime.morestack_noctxt   0�   "".autotmp_0232 �"type.interface {} "".autotmp_0231 �(type.[1]interface {} "".autotmp_0228 /&type.[]interface {} "".autotmp_0227 �type.uint32 "".autotmp_0225 otype."".Value "".autotmp_0224 Otype.string "".autotmp_0223  type.bool "".x �type."".Value "".x �$type."".unknownVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".intVal "".x � type."".int64Val "".~r2 (type.bool "".~r1  type.float32 "".x  type."".Value H����~�����g���� � L�/�O
&�U1LU
5 6 Xsl�p@.Sa�a Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 Tgclocals·82e7e0e6288447ba602a0db7dfa00c79   @$GOROOT/src/go/constant/value.go�"".Float64Val  �  �dH�%    H�D$�H;A�K  H���   W�D$HD$PW�H��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$���T�b  �L$<��1��u~1�H�\$XH�    H�$H��$�   H�\$H��$�   H�\$H�\$XH�\$�    �L$<�\$ �� t5H�\$XH�$�    �D$�\$��$�   �� ��$�   H���   Á��TuzH�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �\$ �� t3H�\$@�H*���$�   �H,�H��H�l$@H9���$�   H���   �H��$�   H��$�   1�H��$�   H��$�   H��$�   H�� �  HǄ$�      HǄ$�      H��$�   H�T$`H�$H�L$hH�L$�    H�L$H�D$H��$�   H�L$pH�H�D$x�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<����>uz1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �L$<�\$ �� t1H�\$HH�$�    �D$�\$��$�   ��$�   H���   Á��|~?u`1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tW���$�   Ƅ$�    H���   Á�@��q�����1�H�\$PH�    H�$H��$�   H�\$H��$�   H�\$H�\$PH�\$�    �\$ �� �g����    H�$H�$H�\$PH�\$�    H�\$H�$�    �D$�\$��$�   �� ��$�   H���   ��    �������4
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  2math/big.(*Float).Float64   �   type."".int64Val   �  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  4go.string."%v not a Float"   �	  fmt.Sprintf   �	  type.string   �
  runtime.convT2E   �
  runtime.gopanic   �
  .runtime.writebarrierptr   �  type."".ratVal   �  $runtime.assertI2T2   �  .math/big.(*Rat).Float64   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  "".newFloat   �  0math/big.(*Float).SetInt   �  2math/big.(*Float).Float64   �  0runtime.morestack_noctxt   @�   "".autotmp_0245 �"type.interface {} "".autotmp_0244 �(type.[1]interface {} "".autotmp_0241 /&type.[]interface {} "".autotmp_0240 �type.uint32 "".autotmp_0238 otype."".Value "".autotmp_0237 Otype.string "".autotmp_0236  type.bool "".x �type."".Value "".x �$type."".unknownVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".intVal "".x � type."".int64Val "".~r2 0type.bool "".~r1  type.float64 "".x  type."".Value J����������g���� � L�/�O
)�U1LU
5 6 Xsl�p@.Sa�^ Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·82e7e0e6288447ba602a0db7dfa00c79   @$GOROOT/src/go/constant/value.go�"".BitLen  �  �dH�%    H�D$�H;A��  H���   1�H�D$HH��$�   H��$�   H��$�   H�$H��$�   H�D$�    �L$�L$<���T��   H�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �L$<�\$ �� t6H�\$@H�$�    H�D$H�D$PH�$�    H�\$H��$�   H���   Á��|~?uX1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tHǄ$�       H���   Á�@��quh1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �\$ �� t#H�\$HH�$�    H�\$H��$�   H���   �H��$�   H��$�   1�H�\$xH��$�   H�\$xH�� �  HǄ$�      HǄ$�      H��$�   H�T$XH�$H�L$`H�L$�    H�L$H�D$H��$�   H�L$hH�H�D$p�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    ������������������(
      �  $runtime.ifacethash   �   type."".int64Val   �  $runtime.assertI2T2   �  "".i64toi   �  ,math/big.(*Int).BitLen   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  ,math/big.(*Int).BitLen   �  runtime.convI2E   �	 (runtime.writeBarrier   �	  2go.string."%v not an Int"   �
  fmt.Sprintf   �
  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   0�  "".autotmp_0257 �"type.interface {} "".autotmp_0256 �(type.[1]interface {} "".autotmp_0253 /&type.[]interface {} "".autotmp_0252 �type.uint32 "".autotmp_0250 otype."".Value "".autotmp_0249 Otype.string "".autotmp_0248  type.int "".autotmp_0246 �type."".intVal "".x �type."".Value "".x �$type."".unknownVal "".x �type."".intVal "".x � type."".int64Val "".~r1  type.int "".x  type."".Value :����_��o���� � 0�&�6LM#� & Omf}{p@.( Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 Tgclocals·9df74eb5f212c312a79ae7ef34903c32   @$GOROOT/src/go/constant/value.go�"".Sign  �  �dH�%    H�D$�H;A�:  H���   W��$�   �$�   D$PD$XH��$�   H��$   H��$�   H�$H��$�   H�D$�    �L$����>�  �L$<��1��ul1�H�\$XH�    H�$H��$�   H�\$H��$�   H�\$H�\$XH�\$�    �L$<�\$ �� t#H�\$XH�$�    H�\$H��$  H���   Á��T��   H�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �L$<�\$ �� tRH�\$@H�� }HǄ$  ����H���   �H�\$@H�� ~HǄ$     H���   �HǄ$      H���   Á���>��   1�H�\$PH�    H�$H��$�   H�\$H��$�   H�\$H�\$PH�\$�    �\$ �� tEH�D$PH�� t6H�hH�� u1�H��$  H���   ���� t	H��������H��   �։ ��H��$�   H��$�   1�H��$�   H��$�   H��$�   H�� �  HǄ$�      HǄ$�      H��$�   H�T$hH�$H�L$pH�L$�    H�L$H�D$H��$�   H�L$xH�H��$�   �=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<���|~?uX1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �L$<�\$ �� tHǄ$     H���   Á�@��q��   1�H�\$`H�    H�$H��$�   H�\$H��$�   H�\$H�\$`H�\$�    �L$<�\$ �� t;H�D$`H�hH�� u1�H��$  H���   ���� t	H��������H��   �ց��q�������1�H��$�   H��$�   H��$�   H��$�   H�    H�$H��$�   H�\$H��$�   H�\$H��$�   H�\$�    �\$ �� �@���H��$�   H�H�$H�KH�L$�    H�\$H�\$HH��$�   H�H�$H�KH�L$�    H�D$H�\$HH	�H��$  H���   ��    ��������4
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  ,math/big.(*Float).Sign   �   type."".int64Val   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �
  runtime.convI2E   � (runtime.writeBarrier   �  4go.string."%v not numeric"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  "".Sign   �  "".Sign   �  0runtime.morestack_noctxt   0�  ("".autotmp_0272 �"type.interface {} "".autotmp_0271 �(type.[1]interface {} "".autotmp_0268 o&type.[]interface {} "".autotmp_0267  type.int "".autotmp_0266 �type.uint32 "".autotmp_0264 �type."".Value "".autotmp_0263 �type.string "".autotmp_0261  type.int "".autotmp_0260  type.int "".autotmp_0259  type.int "".autotmp_0258 �type.int "".x �type."".Value "".x �$type."".unknownVal "".x ?$type."".complexVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".intVal "".x � type."".int64Val "".~r1  type.int "".x  type."".Value l����u������w�����u���� �
 X�<�#WQE�'P$#U;s a! . es^�s@.N�W Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 Tgclocals·8efb4299ccfc450a63c2e51c4c5be655   @$GOROOT/src/go/constant/value.go�"".Bytes  �  �dH�%    H��$x���H;A��  H��  1�H�D$H1�H��$   H��$(  H��$0  1�H�\$PH��$  H��$  H��$�   H�$H��$�   H�D$�    �L$�L$<���T��  H�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �L$<�\$ �� �c  H�\$@H�$�    H�D$H�D$P1�H�� �8  H�hH�XH�HH��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��H��H�    H�$H�D$H�D$�    H�|$L�T$ L�d$(1�H��$�   L��$�   H��$�   E1�M9�}2H�1�H��}L9�s{H��H��H��H��H��|�H��I��M9�|�H�� ~ H��H��L9�sAH�/��� u	H��H�� �L9�w H��$   H��$(  L��$0  H��  ��    �    �    � �������@��quO1�H�\$HH�    H�$H��$�   H�\$H��$�   H�\$H�\$HH�\$�    �\$ �� t
H�D$H�Y���H��$�   H��$�   1�H�\$xH��$�   H�\$xH�� �  HǄ$�      HǄ$      H��$�   H�T$XH�$H�L$`H�L$�    H�L$H�D$H��$�   H�L$hH�H�D$p�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������    �����*
      �  $runtime.ifacethash   �   type."".int64Val   �  $runtime.assertI2T2   �  "".i64toi   �  type.[]uint8   �  "runtime.makeslice   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �	  type."".intVal   �	  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  2go.string."%v not an Int"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   P�  *"".autotmp_0292  type.int "".autotmp_0291  type.int "".autotmp_0289 _(type.[]math/big.Word "".autotmp_0288 �"type.interface {} "".autotmp_0287 �(type.[1]interface {} "".autotmp_0284 /&type.[]interface {} "".autotmp_0283 �type.uint32 "".autotmp_0281 �type."".Value "".autotmp_0279  type.int "".autotmp_0277  type.int "".autotmp_0276  $type.math/big.Word "".autotmp_0275  (type.[]math/big.Word "".autotmp_0273 �type.string "".~r0 �(type.[]math/big.Word "".words �(type.[]math/big.Word "".x �type."".Value "".x �type."".intVal "".x � type."".int64Val "".t �type."".intVal "".~r1  type.[]uint8 "".x  type."".Value ""������ � t�C�]8#	,M
� . sq��Zzp@. Tgclocals·47e744d05637aa546b45723fe9d2d977 Tgclocals·305e11413380417cd9c7d2ae9b79dbaa   @$GOROOT/src/go/constant/value.go� "".MakeFromBytes  �  �dH�%    H;a��  H��h1�H��$�   H��$�   H�\$xH��H��H��?H��=H�H��H��H�    H�$H�D$H�D$�    L�\$L�\$8L�T$ H�\$(H�\$H1�1�1�H�|$pL�d$xH��$�   E1�M9�}R�/I��H��A��H��H��@�,  H��H��H	�H��H��H��@uL9��  I��H�3H��1�1�H��I��M9�|�L�T$@L9���   L9���   I��H�3H��H�D$0H�� ~*H��H��L9���   I��H�H�� uH��H�D$0H�� �H�    H�$�    H�D$H�\$0H�l$HH9�wYL�D$8H�$L�D$PL�D$H�\$XH�\$H�l$`H�l$�    H�\$ H�$�    H�L$H�D$H��$�   H��$�   H��h��    �    �    �4����    1�������    �������������������
      �  (type.[]math/big.Word   �  "runtime.makeslice   �  "type.math/big.Int   �  "runtime.newobject   �  .math/big.(*Int).SetBits   �  "".makeInt   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   P�  "".autotmp_0310  type.int "".autotmp_0309  type.int "".autotmp_0307  type.int "".autotmp_0305  $type.*math/big.Int "".autotmp_0304 /(type.[]math/big.Word "".autotmp_0302  type.int "".autotmp_0301  type.int "".autotmp_0300  type.int "".i otype.int "".words _(type.[]math/big.Word "".~r1 0type."".Value "".bytes  type.[]uint8  ����(� � n�)Q  
'�  \�@s Tgclocals·3260b5c802f633fd6252c227878dd72a Tgclocals·524aafe7d1228e5424d64f5d94771fbf   @$GOROOT/src/go/constant/value.go�"".Num  �  �dH�%    H�D$�H;A�c  H��   W�D$@1�H��$�   H��$�   H��$�   H��$�   H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �L$���T��  �L$<��1���  1�H�\$HH�    H�$H�T$H�l$H�\$HH�\$�    H��$�   H��$�   �L$<�\$ �� ��   H�\$HH�$�    �\$�� tQH�\$HH�$H�D$    �    H�\$H�� t+H�$�    H�L$H�D$H��$�   H��$�   H�ĸ   É��1�H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�   H�\$0H��$�   H�ĸ   Á��TuUH�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �\$ �� tH��$�   H��$�   H�ĸ   �1�H�\$pH�\$xH�\$pH�� �  HǄ$�      HǄ$�      H��$�   H�T$PH�$H�l$XH�l$�    H�L$H�D$H��$�   H�L$`H�H�D$h�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<����>��   1�H�\$@H�    H�$H�T$H�l$H�\$@H�\$�    H��$�   H��$�   �L$<�\$ �� t:H�\$@H�� t+H�$�    H�L$H�D$H��$�   H��$�   H�ĸ   É�с��|~?uH1�H�    H�$H�T$H�l$H�\$<H�\$�    H��$�   H��$�   �L$<�\$ �� �$�����@��q�����H�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �\$ �� �{��������    �{��������������:
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  "".smallRat   �  *math/big.(*Float).Rat   �  "".makeInt   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �   type."".int64Val   �  $runtime.assertI2T2   �	  runtime.convI2E   �	 (runtime.writeBarrier   �
  >go.string."%v not Int or Float"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  type."".ratVal   �  $runtime.assertI2T2   �  "".makeInt   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   @�   "".autotmp_0327 �"type.interface {} "".autotmp_0326 �(type.[1]interface {} "".autotmp_0323 /&type.[]interface {} "".autotmp_0322  $type.*math/big.Int "".autotmp_0320 �type.uint32 "".autotmp_0318 otype."".Value "".autotmp_0317 �$type."".unknownVal "".autotmp_0316 Otype.string "".autotmp_0315  type."".Value "".autotmp_0314  type.bool "".x �type."".Value "".x �$type."".unknownVal "".x � type."".floatVal "".x �type."".ratVal "".~r1  type."".Value "".x  type."".Value H����b��\������� �	 B�	9�5_E�Y:� 6 b���p@.G2T� Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·0000613cea0d43cb0624ba62b8fe2aca   @$GOROOT/src/go/constant/value.go�"".Denom  �  �dH�%    H�D$�H;A��  H���   W�D$H1�H��$�   H��$�   H��$�   H��$�   H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �L$���T�+  �L$<��1���  1�H�\$PH�    H�$H�T$H�l$H�\$PH�\$�    H��$�   H��$�   �L$<�\$ �� ��   H�\$PH�$�    �\$�� tUH�\$PH�$H�D$    �    H�\$H�$�    H�\$H�$�    H�L$H�D$H��$�   H��$�   H���   �1�H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�   H�\$0H��$�   H���   Á��T��   H�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �\$ �� tpH�T$XH�l$`H�D$@   H�    H�$H�    H�\$H�    H�\$H�\$@H�\$H�D$     �    H�\$(H��$�   H�\$0H��$�   H���   �1�H��$�   H��$�   H��$�   H�� �  HǄ$�      HǄ$�      H��$�   H�T$hH�$H�l$pH�l$�    H�L$H�D$H��$�   H�L$xH�H��$�   �=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<����>��   1�H�\$HH�    H�$H�T$H�l$H�\$HH�\$�    H��$�   H��$�   �L$<�\$ �� t>H�\$HH�$�    H�\$H�$�    H�L$H�D$H��$�   H��$�   H���   Á��|~?uH1�H�    H�$H�T$H�l$H�\$<H�\$�    H��$�   H��$�   �L$<�\$ �� �������@��q�����H�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �\$ �� �����~����    ���������������F
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  "".smallRat   �  *math/big.(*Float).Rat   �  *math/big.(*Rat).Denom   �  "".makeInt   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �   type."".int64Val   �  $runtime.assertI2T2   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �	  runtime.convT2I   �  runtime.convI2E   � (runtime.writeBarrier   �  >go.string."%v not Int or Float"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  type."".ratVal   �  $runtime.assertI2T2   �  *math/big.(*Rat).Denom   �  "".makeInt   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   @�  $"".autotmp_0343 �"type.interface {} "".autotmp_0342 �(type.[1]interface {} "".autotmp_0339 /&type.[]interface {} "".autotmp_0338 �type.uint32 "".autotmp_0336 otype."".Value "".autotmp_0335 �$type."".unknownVal "".autotmp_0334 Otype.string "".autotmp_0333  type."".Value "".autotmp_0332  $type.*math/big.Int "".autotmp_0331  type.bool "".autotmp_0328 � type."".int64Val "".x �type."".Value "".x �$type."".unknownVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".Value "".~r1  type."".Value "".x  type."".Value J����^���������� �
 F�	9�9_I
f�Y>� 8 b��h~s@.G,^� Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·c04ada1956856a77e3bc187a9e8a1dcc   @$GOROOT/src/go/constant/value.go�"".MakeImag  �  �dH�%    H�D$�H;A�x  H���   1�H��$  H��$  H��$�   H��$   H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �L$���T�  �L$<��1���u  H�    H�$H�l$H�T$H�D$    �    H��$�   H��$�   �L$<�\$ �� �0  H�D$@    H�    H�$H�    H�\$H�    H�\$H�\$@H�\$H�D$     �    H�l$(H�T$0H��$�   H��$�   H��$�   H��$   1�H�\$HH�\$P1�H��$�   H��$�   H��$�   H��$�   H�l$XH��$�   H�T$`H��$�   H�L$hH��$�   H�D$pH��$�   H�    H�$H�    H�\$H�    H�\$H��$�   H�\$H�D$     �    H�L$(H�D$0H��$  H��$  H���   Á��Tu1H�    H�$H�l$H�T$H�D$    �    �\$ �� �����1�H��$�   H��$�   H��$�   H�� �$  HǄ$�      HǄ$�      H��$�   H��$�   H�$H��$   H�\$�    H�L$H�D$H��$�   H�L$xH�H��$�   �=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<����>uEH�    H�$H�l$H�T$H�D$    �    H��$�   H��$�   �L$<�\$ �� ��������|~?uiH�    H�$H�l$H�T$H�D$    �    H��$�   H��$�   �L$<�\$ �� t(H��$�   H��$  H��$   H��$  H���   Á�@��q�����H�    H�$H�l$H�T$H�D$    �    �\$ �� �I��������    �f���������:
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �   type."".int64Val   �  $runtime.assertI2T2   �
  runtime.convI2E   � (runtime.writeBarrier   �  >go.string."%v not Int or Float"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  type."".ratVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   @�  "".autotmp_0356 �"type.interface {} "".autotmp_0355 �(type.[1]interface {} "".autotmp_0352 o&type.[]interface {} "".autotmp_0351  type."".Value "".autotmp_0350  type."".Value "".autotmp_0349 �type.uint32 "".autotmp_0347 �type."".Value "".autotmp_0346 �type.string "".autotmp_0345 ?$type."".complexVal "".autotmp_0344 � type."".int64Val "".~r2 �type."".Value 
"".im �type."".Value 
"".re �type."".Value "".~r1  type."".Value "".x  type."".Value .�������B� �	 4�	1��9��(= 4 Z��Mps@.;�( Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·5ff70dccce69b73e733742f8f6b97bd8   @$GOROOT/src/go/constant/value.go�"".Real  �  �dH�%    H�D$�H;A��  H���   W��$�   �$�   1�H��$�   H��$�   H��$�   H��$�   H�L$pH�$H�D$xH�D$�    H�T$pH�l$x�L$����>�"  �L$<��1��uSH�    H�$H�T$H�l$H�D$    �    H�T$pH�l$x�L$<�\$ �� tH��$�   H��$�   H���   Á��Tu;H�    H�$H�T$H�l$H�D$    �    H�T$pH�l$x�L$<�\$ �� u�����>u;H�    H�$H�T$H�l$H�D$    �    H�T$pH�l$x�\$ �� �b���1�H�\$`H�\$hH�\$`H�� �  HǄ$�      HǄ$�      H��$�   H�T$@H�$H�l$HH�l$�    H�L$H�D$H��$�   H�L$PH�H�D$X�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<���|~?u?H�    H�$H�T$H�l$H�D$    �    H�T$pH�l$x�L$<�\$ �� �������@��qu?H�    H�$H�T$H�l$H�D$    �    H�T$pH�l$x�L$<�\$ �� ��������q���%���1�H��$�   H��$�   H��$�   H��$�   H�    H�$H�T$H�l$H��$�   H�\$�    H�T$pH�l$x�\$ �� �����H��$�   H��$�   H��$�   H��$�   H���   ��    �'����������.
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �  runtime.convI2E   � (runtime.writeBarrier   �  4go.string."%v not numeric"   �  fmt.Sprintf   �	  type.string   �	  runtime.convT2E   �
  runtime.gopanic   �
  .runtime.writebarrierptr   �
  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   @�  "".autotmp_0365 �"type.interface {} "".autotmp_0364 �(type.[1]interface {} "".autotmp_0361 o&type.[]interface {} "".autotmp_0360 �type.uint32 "".autotmp_0358 �type."".Value "".autotmp_0357 �type.string "".x �type."".Value "".x ?$type."".complexVal "".~r1  type."".Value "".x  type."".Value "������ � ,�
D����(	 " g�p@.;� Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc Tgclocals·2bee6dd56e8b158e514a8950bd21767b   @$GOROOT/src/go/constant/value.go�"".Imag  �  �dH�%    H�D$�H;A��  H���   W��$�   �$�   1�H��$�   H��$   H��$�   H��$�   H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �L$����>��  �L$<��1����   H�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �L$<�\$ �� tpH�T$XH�l$`H�D$@    H�    H�$H�    H�\$H�    H�\$H�\$@H�\$H�D$     �    H�\$(H��$�   H�\$0H��$   H���   Á��TuEH�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �L$<�\$ �� �C�������>uAH�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �\$ �� �����1�H�\$xH��$�   H�\$xH�� �  HǄ$�      HǄ$�      H��$�   H�T$HH�$H�l$PH�l$�    H�L$H�D$H��$�   H�L$hH�H�D$p�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M����������L$<���|~?��   1�H�    H�$H�T$H�l$H�\$<H�\$�    H��$�   H��$�   �L$<�\$ �� t]H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�   H�\$0H��$   H���   Á�@��quEH�    H�$H�T$H�l$H�D$    �    H��$�   H��$�   �L$<�\$ �� ��������q�������1�H��$�   H��$�   H��$�   H��$�   H�    H�$H�T$H�l$H��$�   H�\$�    H��$�   H��$�   �\$ �� �O���H��$�   H��$�   H��$�   H��$   H���   ��    �4�������>
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �   type."".int64Val   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �  runtime.convI2E   �	 (runtime.writeBarrier   �	  4go.string."%v not numeric"   �
  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  $type."".unknownVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  type."".intVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   @�  "".autotmp_0376 �"type.interface {} "".autotmp_0375 �(type.[1]interface {} "".autotmp_0372 o&type.[]interface {} "".autotmp_0371 �type.uint32 "".autotmp_0369 �type."".Value "".autotmp_0368 �type.string "".autotmp_0367 � type."".int64Val "".autotmp_0366 �$type."".unknownVal "".x �type."".Value "".x ?$type."".complexVal "".x �type."".Value "".x �$type."".unknownVal "".~r1  type."".Value "".x  type."".Value 0��������� �	 8�
D�
f��T]�( 4 m�M�p@.BYM� Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·707962cf7cb527a8361df5d978b0d876   @$GOROOT/src/go/constant/value.go�"".ToInt  �  �dH�%    H�D$�H;A��  H���   W��$�   �$�   �$�   D$x�$�   D$@1�H��$�   H��$   H��$�   H��$�   H�L$hH�$H�D$pH�D$�    H�l$hH�T$p�L$���T��  �L$<��1���g  1�H�\$@H�    H�$H�l$H�T$H�\$@H�\$�    H�l$hH�T$p�L$<�\$ �� �   H�\$@H�$�    �\$�� �  H�    H�$�    H�D$H�\$@H�$H�D$PH�D$�    �\$�� u0H�\$PH�$�    H�L$H�D$H��$�   H��$   H���   �H��$�   W�CCH��$�   H�$H�D$�  �    H��$�   H��   �K�C H��$�   H�$H�\$@H�\$�    H��$�   H�$H�\$PH�\$�    �\$�� u0H�\$PH�$�    H�L$H�D$H��$�   H��$   H���   �H��$�   H��   �K�C H��$�   H�$H�\$@H�\$�    H��$�   H�$H�\$PH�\$�    �\$�� u0H�\$PH�$�    H�L$H�D$H��$�   H��$   H���   �1�H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�   H�\$0H��$   H���   �럁��Tu�H�    H�$H�l$H�T$H�D$    �    H�l$hH�T$p�\$ �� �\���H��$�   H��$   H���   ÉL$<����>��   1�H�\$HH�    H�$H�l$H�T$H�\$HH�\$�    H�l$hH�T$p�L$<�\$ �� tWH�\$HH�$�    �\$�� t:H�\$HH�� t+H�$�    H�L$H�D$H��$�   H��$   H���   É��������@��qu?H�    H�$H�l$H�T$H�D$    �    H�l$hH�T$p�L$<�\$ �� ��������q���G���1�H�\$xH��$�   H��$�   H��$�   H�    H�$H�l$H�T$H�\$xH�\$�    �\$ �� �����H�\$xH��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H�    H�$H�    H�\$H�    H�\$H��$�   H�\$H�D$     �    H�\$(H�H�$H�KH�L$�    H�L$H�D$H�D$`H�$H�L$XH�Y(��H�\$H��u:H�\$XH�$H�\$`H�\$�    H�L$H�D$H��$�   H��$   H���   �������    �9������������L
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  "".smallRat   �  "type.math/big.Int   �  "runtime.newobject   �  *math/big.(*Float).Int   �  "".makeInt   �  2math/big.(*Float).SetPrec   �  *math/big.(*Float).Set   �  *math/big.(*Float).Int   �  "".makeInt   �	  *math/big.(*Float).Set   �	  *math/big.(*Float).Int   �
  "".makeInt   �
  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �   type."".int64Val   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �  *math/big.(*Rat).IsInt   �  "".makeInt   �  type."".intVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �  "".ToFloat   �       �  "".ToInt   �  0runtime.morestack_noctxt   @�  ("".autotmp_0390 �type.uint32 "".autotmp_0388 �type."".Value "".autotmp_0387 �$type."".unknownVal "".autotmp_0386  type."".Value "".autotmp_0384 �$type."".complexVal "".autotmp_0383  type."".Value "".autotmp_0382  type."".Value "".autotmp_0381  type."".Value "".autotmp_0380  $type.*math/big.Int "".autotmp_0379  type.bool "".autotmp_0378  type."".Value "".autotmp_0377  type.bool 
"".re �type."".Value "".x �$type."".complexVal "".t O&type.math/big.Float "".i �$type.*math/big.Int "".x � type."".floatVal "".x �type."".ratVal "".~r1  type."".Value "".x  type."".Value p����������^��\��������� � z�
^�"0%0%0a_CS
:T_�V�:a J �;RdS3��tk�; ? Tgclocals·a68b09a48716afad7ca7a02fe6add474 Tgclocals·5a22249a9b0f12f04d737839c0e5b8d8   @$GOROOT/src/go/constant/value.go�"".ToFloat  �  �dH�%    H�D$�H;A��  H��   W�D$x�$�   1�H�D$H1�H��$�   H��$�   H��$�   H��$�   H�L$hH�$H�D$pH�D$�    H�l$hH�T$p�L$���T�s  �L$<��1��uSH�    H�$H�l$H�T$H�D$    �    H�l$hH�T$p�L$<�\$ �� tH��$�   H��$�   H�Ę   Á��T��   H�D$@    H�    H�$H�l$H�T$H�\$@H�\$�    �\$ �� trH�\$@H�$�    H�\$H�\$PH�    1�H9�tH�\$PH��$�   H��$�   H�Ę   �H�    H�$H�    H�\$H�    H�\$�    H�D$�1�H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�   H�\$0H��$�   H�Ę   ÉL$<����>u?H�    H�$H�l$H�T$H�D$    �    H�l$hH�T$p�L$<�\$ �� �������@��q��   1�H�\$HH�    H�$H�l$H�T$H�\$HH�\$�    H�l$hH�T$p�L$<�\$ �� trH�\$HH�$�    H�\$H�\$PH�    1�H9�tH�\$PH��$�   H��$�   H�Ę   �H�    H�$H�    H�\$H�    H�\$�    H�D$봁��q�������1�H�\$xH��$�   H��$�   H��$�   H�    H�$H�l$H�T$H�\$xH�\$�    �\$ �� �8���H��$�   H�H�$H�KH�L$�    H�L$H�D$H�D$`H�$H�L$XH�Y(��H�\$H��u_H�\$XH�$H�\$`H�\$�    H�\$H�� u<H�\$xH�H�$H�KH�L$�    H�L$H�D$H��$�   H��$�   H�Ę   ������    �����������B
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  $runtime.assertI2T2   �  "".i64tof   �  8go.itab."".floatVal."".Value   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  type."".ratVal   �  $runtime.assertI2T2   �	  type."".intVal   �	  $runtime.assertI2T2   �
  "".itof   �
  8go.itab."".floatVal."".Value   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  $type."".complexVal   �  $runtime.assertI2T2   �  "".ToInt   �       �  "".Sign   �  "".ToFloat   �  0runtime.morestack_noctxt   @�  "".autotmp_0402  type.*uint8 "".autotmp_0400 �type.uint32 "".autotmp_0398 _type."".Value "".autotmp_0397 �$type."".unknownVal "".autotmp_0396  type."".Value "".autotmp_0393   type."".floatVal "".autotmp_0392 � type."".floatVal 
"".im type."".Value "".x ?$type."".complexVal "".x �type."".intVal "".x � type."".int64Val "".~r1  type."".Value "".x  type."".Value X����������������� � <�H�Cr_�r]i< 0 k�uDQy]VL a Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc Tgclocals·9d7301afadfdafb7e149f098ce5d5791   @$GOROOT/src/go/constant/value.go�"".ToComplex  �,  �,dH�%    H��$����H;A��
  H��  W��$H  �$X  D$PD$X1�H��$�  H��$�  H��$�  H��$�  H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �L$���T��  �L$<��1���4  1�H�\$XH�    H�$H�l$H�T$H�\$XH�\$�    H��$�   H��$�   �L$<�\$ �� ��  H�\$XH�\$pH�    1�H9���  H�T$pH��$�   H��$�   1�H��$(  H��$0  H��$8  H��$@  H�D$H    1�H��$h  H��$p  H��$x  H��$�  H��$�   H��$h  H��$�   H��$p  H�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�\$(H��$x  H�H�M H�KH�MH��$h  H��$p  H��$x  H��$�  H��$(  H��$�  H��$0  H��$�  H��$8  H��$�  H��$@  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  �H�    H�$H�    H�\$H�    H�\$�    H�D$�5������T�-  H�D$@    H�    H�$H�l$H�T$H�\$@H�\$�    �\$ �� ��  H�\$@H�$�    H�\$H�\$pH�    1�H9���  H�T$pH��$�   H��$�   1�H��$�   H��$�   H��$�   H��$   H�D$H    1�H��$h  H��$p  H��$x  H��$�  H�D$xH��$h  H��$�   H��$p  H�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�\$(H��$x  H�H�M H�KH�MH��$h  H��$p  H��$x  H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H��$   H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  �H�    H�$H�    H�\$H�    H�\$�    H�D$�8���1�H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  ÉL$<����>�4  1�H�\$PH�    H�$H�l$H�T$H�\$PH�\$�    H��$�   H��$�   �L$<�\$ �� ��  H�\$PH�\$hH�    1�H9���  H�T$hH��$�   H��$�   1�H��$  H��$  H��$  H��$   H�D$H    1�H��$h  H��$p  H��$x  H��$�  H��$�   H��$h  H��$�   H��$p  H�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�\$(H��$x  H�H�M H�KH�MH��$h  H��$p  H��$x  H��$�  H��$  H��$�  H��$  H��$�  H��$  H��$�  H��$   H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  �H�    H�$H�    H�\$H�    H�\$�    H�D$�5�����@��q�B  1�H�\$`H�    H�$H�l$H�T$H�\$`H�\$�    H��$�   H��$�   �L$<�\$ �� ��  H�\$`H�$�    H�\$H�\$pH�    1�H9���  H�T$pH��$�   H��$�   1�H��$�   H��$�   H��$�   H��$�   H�D$H    1�H��$h  H��$p  H��$x  H��$�  H��$�   H��$h  H��$�   H��$p  H�    H�$H�    H�\$H�    H�\$H�\$HH�\$H�D$     �    H�\$(H��$x  H�H�M H�KH�MH��$h  H��$p  H��$x  H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  �H�    H�$H�    H�\$H�    H�\$�    H�D$�5������q������1�H��$H  H��$P  H��$X  H��$`  H�    H�$H�l$H�T$H��$H  H�\$�    �\$ �� �����H��$H  H��$�  H��$P  H��$�  H��$X  H��$�  H��$`  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H�Ĩ  ��    ����������̖
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  8go.itab."".floatVal."".Value   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �	  $type."".complexVal   �	  type."".Value   �	  <go.itab."".complexVal."".Value   �
  runtime.convT2I   �
   type."".floatVal   �
  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �   type."".int64Val   �  $runtime.assertI2T2   �  "".i64tof   �  8go.itab."".floatVal."".Value   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  type."".ratVal   �  $runtime.assertI2T2   �  4go.itab."".ratVal."".Value   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �  type."".ratVal   �  type."".Value   �  4go.itab."".ratVal."".Value   �   runtime.typ2Itab   �  type."".intVal   �  $runtime.assertI2T2   �   "".itof   �   8go.itab."".floatVal."".Value   �#   type."".int64Val   �#  type."".Value   �#  8go.itab."".int64Val."".Value   �#  runtime.convT2I   �%  $type."".complexVal   �&  type."".Value   �&  <go.itab."".complexVal."".Value   �&  runtime.convT2I   �'   type."".floatVal   �'  type."".Value   �'  8go.itab."".floatVal."".Value   �'   runtime.typ2Itab   �(  $type."".complexVal   �)  $runtime.assertI2T2   �*  $type."".complexVal   �*  type."".Value   �+  <go.itab."".complexVal."".Value   �+  runtime.convT2I   �,  0runtime.morestack_noctxt   @�  T"".autotmp_0433  $type."".complexVal "".autotmp_0432  type.*uint8 "".autotmp_0431  type."".Value "".autotmp_0430  $type."".complexVal "".autotmp_0429  type.*uint8 "".autotmp_0428  type."".Value "".autotmp_0427  $type."".complexVal "".autotmp_0426  type.*uint8 "".autotmp_0425  type."".Value "".autotmp_0424 $type."".complexVal "".autotmp_0422  type."".Value "".autotmp_0421 �type.uint32 "".autotmp_0419 �type."".Value "".autotmp_0418 �$type."".unknownVal "".autotmp_0417  $type."".complexVal "".autotmp_0416  $type."".complexVal "".autotmp_0415   type."".int64Val "".autotmp_0414   type."".floatVal "".autotmp_0413  $type."".complexVal "".autotmp_0412   type."".int64Val "".autotmp_0411 �type."".ratVal "".autotmp_0410  $type."".complexVal "".autotmp_0409   type."".int64Val "".autotmp_0408   type."".floatVal "".autotmp_0407 ?$type."".complexVal "".autotmp_0406 � type."".int64Val "".autotmp_0405 � type."".floatVal "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".x �$type."".complexVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".intVal "".x � type."".int64Val "".~r1  type."".Value "".x  type."".Value Z"������������������ � D�Q��G�_]�Y�c� h z��JC��JG]��JA	0��J_�7 Tgclocals·1dbe3e1675327063a63a3ea108cf04bf Tgclocals·ba07643250a35734cb355a9fec6f55cc   @$GOROOT/src/go/constant/value.go�"".is32bit  @  @H�D$H=   �|H=����D$��D$ ��     "".~r1 type.bool "".x  type.int64     �  Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".is63bit  `  `H�D$H�       �H9�|H��������?H9��D$��D$ ����     "".~r1 type.bool "".x  type.int64 0 0 �+  Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".UnaryOp  �<  �<dH�%    H��$����H;A��  H���  W��$�  �$�  �$@  �$P  D$x�$�   H��$�  H��$�  1�H��$�  H��$�  H��$�  H���
  H����  H��$  H�$H��$  H�L$�    H��$  H��$  �L$����>��  �L$<��1��uiH�    H�$H�l$H�T$H�D$    �    H��$  H��$  �L$<�\$ �� t(H��$�  H��$�  H��$�  H��$�  H���  Á��TuAH�    H�$H�l$H�T$H�D$    �    H��$  H��$  �L$<�\$ �� u�����>u1H�    H�$H�l$H�T$H�D$    �    �\$ �� �V���H��$�  H�\$P1�H��$`  H��$h  H��$p  H��$x  H��$`  H�� ��  HǄ$0     HǄ$8     H��$(  H�    H�$H�\$PH�\$H�D$    �    H�L$H�D$ H��$(  H��$�   H�H��$   �=     �  H�CH��$�  H�$H��$�  H�\$�    H�L$H�D$H��$(  H��H��$�   H�H��$   �=     ��   H�CH�    H�$H�D$   H��$(  H�\$H��$0  H�\$H��$8  H�\$ �    H�\$(H��$  H�\$0H��$   H�    H�$H��$  H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M���L�CL�$H�D$�    �������^����L$<���|~?uEH�    H�$H�l$H�T$H�D$    �    H��$  H��$  �L$<�\$ �� �"�����@��quEH�    H�$H�l$H�T$H�D$    �    H��$  H��$  �L$<�\$ �� ��������q���s���H�    H�$H�l$H�T$H�D$    �    �\$ �� ������=���H���3���H��$  H�$H��$  H�L$�    H��$  H��$  �L$����>��  �L$<��1����   1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$  H��$  �L$<�\$ �� tO�    H�$H�$H��$�   H�\$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H���  Á��T�3  H�D$H    H�    H�$H�l$H�T$H�\$HH�\$�    H��$  H��$  �L$<�\$ �� ��   H�D$HH��H�l$HH9�tbH�D$XH�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H���  �H�    H�$�    H�\$H�\$`H�\$HH�$�    H�D$H�\$`H�$H�D$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H���  Á���>�����1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    �\$ �� �����H�    H�$�    H�\$H�$H��$�   H�\$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H���  ÉL$<���|~?��   1�H�    H�$H�l$H�T$H�\$:H�\$�    H��$  H��$  �L$<�\$ �� t]H�    H�$H�    H�\$H�    H�\$H�\$:H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H���  Á�@��q��   1�H�\$xH�    H�$H�l$H�T$H�\$xH�\$�    H��$  H��$  �L$<�\$ �� tXH�    H�$�    H�\$H�$H�\$xH�\$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H���  Á��q�������1�H��$@  H��$H  H��$P  H��$X  H�    H�$H�l$H�T$H��$@  H�\$�    �\$ �� �����H�$   H��$@  H�|$H�H�H�KH�OH�D$    �    H�\$ H��$�   H�\$(H��$�   H�$   H��$P  H�|$H�H�H�KH�OH�D$    �    H�L$ H�D$(H��$�   H��$�   H��$�   H��$�   1�H��$�   H��$�   1�H��$�  H��$�  H��$�  H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H��$�   H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$�  H��$�  H���  �H����  H�    H�$�    H�\$H�\$pH��$�  H��$�  H��$  H�$H��$  H�D$�    �L$�L$<���T�0  H�D$@    H�    H�$H��$  H�\$H��$  H�\$H�\$@H�\$�    �L$<�\$ �� ��   H�\$@H�$�    H�D$H�\$pH�$H�D$�    H��$�  H�� v}1ۈ�$�  H��$�  H��$�  H��$�  H��$�  H�\$hH�$�����    H�D$H�\$hH�$H�D$H��$�  H�\$�    H�L$pH�D$H�$H�L$H�D$�    H�\$pH�$�    H�L$H�D$H��$�  H��$�  H���  Á��|~?��   1�H�    H�$H��$  H�\$H��$  H�\$H�\$:H�\$�    �L$<�\$ �� t]H�    H�$H�    H�\$H�    H�\$H�\$:H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H���  Á�@��quk1�H��$�   H�    H�$H��$  H�\$H��$  H�\$H��$�   H�\$�    �\$ �� t H�\$pH�$H��$�   H�\$�    �%���H��$  H��$�   H��$  H��$�   �L���H��+�B���H��$  H�$H��$  H�L$�    �L$�L$<����
&��   �D$: H�    H�$H��$  H�\$H��$  H�\$H�\$:H�\$�    �L$<�\$ �� tk�\$:�\$;�t$;H�    H�$H�    H�\$H�    H�\$H�\$;H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H���  Á��|~?�R���1�H�    H�$H��$  H�\$H��$  H�\$H�\$:H�\$�    �\$ �� ����H�    H�$H�    H�\$H�    H�\$H�\$:H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H���  ��    ��������
      �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �  &type.go/token.Token   �	  runtime.convT2E   �	 (runtime.writeBarrier   �
  runtime.convI2E   � (runtime.writeBarrier   �  Pgo.string."invalid unary operation %s%v"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  "".newFloat   �  *math/big.(*Float).Neg   �  "".makeFloat   �   type."".int64Val   �  $runtime.assertI2T2   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "type.math/big.Int   �  "runtime.newobject   �  math/big.NewInt   �  &math/big.(*Int).Neg   �  "".makeInt   �  type."".ratVal   �  $runtime.assertI2T2   �  "type.math/big.Rat   �  "runtime.newobject   �  &math/big.(*Rat).Neg   �  "".makeRat   �  $type."".unknownVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �   type."".intVal   �!  $runtime.assertI2T2   �!  "type.math/big.Int   �!  "runtime.newobject   �"  &math/big.(*Int).Neg   �"  "".makeInt   �#  $type."".complexVal   �$  $runtime.assertI2T2   �%  "".UnaryOp   �&  "".UnaryOp   �)  $type."".complexVal   �)  type."".Value   �)  <go.itab."".complexVal."".Value   �)  runtime.convT2I   �*  "type.math/big.Int   �*  "runtime.newobject   �+  $runtime.ifacethash   �,   type."".int64Val   �,  $runtime.assertI2T2   �-  math/big.NewInt   �-  &math/big.(*Int).Not   �.  math/big.NewInt   �/  &math/big.(*Int).Lsh   �0  ,math/big.(*Int).AndNot   �0  "".makeInt   �1  $type."".unknownVal   �1  $runtime.assertI2T2   �2  $type."".unknownVal   �2  type."".Value   �2  <go.itab."".unknownVal."".Value   �2  runtime.convT2I   �3  type."".intVal   �4  $runtime.assertI2T2   �5  &math/big.(*Int).Not   �6  $runtime.ifacethash   �6  type."".boolVal   �7  $runtime.assertI2T2   �8  type."".boolVal   �8  type."".Value   �8  6go.itab."".boolVal."".Value   �9  runtime.convT2I   �9  $type."".unknownVal   �:  $runtime.assertI2T2   �:  $type."".unknownVal   �;  type."".Value   �;  <go.itab."".unknownVal."".Value   �;  runtime.convT2I   �<  0runtime.morestack_noctxt   `�  �"".autotmp_0485  "type.interface {} "".autotmp_0484 �"type.interface {} "".autotmp_0483 �(type.[2]interface {} "".autotmp_0480 �&type.[]interface {} "".autotmp_0479  type.uint32 "".autotmp_0478  type.bool "".autotmp_0477  type."".Value "".autotmp_0476 "type.math/big.Int "".autotmp_0475  type.uint32 "".autotmp_0474  type.bool "".autotmp_0473  type."".Value "".autotmp_0472  type."".Value "".autotmp_0471  type.uint32 "".autotmp_0470  type.bool "".autotmp_0469  type."".Value "".autotmp_0468 �type.uint32 "".autotmp_0466 �type."".Value "".autotmp_0464 �type.string "".autotmp_0463 �&type.go/token.Token "".autotmp_0462 �type."".boolVal "".autotmp_0461  $type."".unknownVal "".autotmp_0460  type."".Value "".autotmp_0458  $type.*math/big.Int "".autotmp_0457  $type.*math/big.Int "".autotmp_0456  $type.*math/big.Int "".autotmp_0455  $type."".unknownVal "".autotmp_0454  $type.*math/big.Int "".autotmp_0453 ?$type."".complexVal "".autotmp_0452  type."".Value "".autotmp_0451  (type.*math/big.Float "".autotmp_0449  type."".Value "".autotmp_0448  $type.*math/big.Rat "".autotmp_0446  type."".Value "".autotmp_0445  $type.*math/big.Int "".autotmp_0444  $type.*math/big.Int "".autotmp_0443  type."".Value "".autotmp_0442  $type.*math/big.Int "".autotmp_0441  $type.*math/big.Int "".autotmp_0439 � type."".int64Val "".autotmp_0438 �$type."".unknownVal "".~r0 �$type.*math/big.Int "".~r2 �type."".Value 
"".im �type."".Value 
"".re �type."".Value "".~r0 �$type.*math/big.Int "".y �type."".boolVal "".y �$type."".unknownVal "".y �type."".Value "".y �type."".intVal "".y � type."".int64Val "".y �$type."".unknownVal "".z �$type.*math/big.Int 
"".im �type."".Value 
"".re �type."".Value "".y �$type."".complexVal "".y � type."".floatVal "".y �type."".ratVal "".y �type."".intVal "".y � type."".int64Val "".y �$type."".unknownVal "".~r3 @type."".Value "".prec 0type.uint "".y type."".Value 
"".op  &type.go/token.Token �"����������o������������������������� � ��t
�(�p�o�pe
�O[bpK[T]UXcK;�
�&}0P]S *
ykP]g � ����@.R�;��tJ�YY.��<8qa%+	dIk%R�� Tgclocals·33962f28c07936e169c43edefa5ca65b Tgclocals·37508b3b9062b4dfe185a1b1456475c6   @$GOROOT/src/go/constant/value.go�"".ord  �  �dH�%    H;a�  H��PH�L$XH�D$`H�L$0H�$H�D$8H�D$�    H�T$0H�L$8�D$=��>��  =�T��   �D$,=1��uIH�    H�$H�T$H�L$H�D$    �    H�T$0H�L$8�D$,�\$ �� tH�D$h   H��P�=�Tu;H�    H�$H�T$H�L$H�D$    �    �\$ �� tH�D$h   H��P�H�    H�\$@H�D$H   H�    H�$H�\$@H�\$H�D$    �    H�\$H�H�$H�KH�L$�    �D$,=��
&uIH�    H�$H�T$H�L$H�D$    �    H�T$0H�L$8�D$,�\$ �� tH�D$h   H��P�=��>�M���H�    H�$H�T$H�L$H�D$    �    �\$ �� ����H�D$h   H��P�=@��q��   �D$,=�|~?uIH�    H�$H�T$H�L$H�D$    �    H�T$0H�L$8�D$,�\$ �� tH�D$h    H��P�=@��q�����H�    H�$H�T$H�L$H�D$    �    �\$ �� �s���H�D$h   H��PÉD$,=�n�u?H�    H�$H�T$H�L$H�D$    �    H�T$0H�L$8�D$,�\$ �� �����=�q������H�    H�$H�T$H�L$H�D$    �    �\$ �� �����H�D$h   H��P��    ���������.
      j  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".int64Val   �  $runtime.assertI2T2   �  .go.string."unreachable"   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  type."".boolVal   �  $runtime.assertI2T2   �  type."".ratVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  $runtime.assertI2T2   �	  type."".intVal   �	  $runtime.assertI2T2   �
  "type."".stringVal   �
  $runtime.assertI2T2   �  $type."".complexVal   �  $runtime.assertI2T2   �  0runtime.morestack_noctxt   0�  
"".autotmp_0489 Gtype.uint32 "".autotmp_0487 ?type."".Value "".autotmp_0486 type.string "".~r1  type.int "".x  type."".Value `����A�����I��^��I���� � L��4TF<Q<� , 4�PJTUTJJ/ Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 Tgclocals·e94709487fd39cb5e22f0477cb3700dd   @$GOROOT/src/go/constant/value.go�"".match  �  �dH�%    H��$����H;A��  H���  W�H��$  �    H�|$P�    1�1�1�H��$(  H��$0  1�H��$  H��$   H��$�  H�$H��$   H�\$�    H�\$H�\$hH��$  H�$H��$  H�\$�    H��$�  H��$   H�D$H�\$hH9�~dH��$  H�$H��$  H�\$H�L$H�T$�    H�L$ H�D$(H�l$0H�T$8H��$  H��$   H��$(  H��$0  H���  �H��$p  H�$H��$x  H�T$�    H��$p  H��$x  �D$=��>��  =�T�$  �D$D=1���M  1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    H��$p  H��$x  �D$D�\$ �� ��  H��$  H��$  H��$P  H�$H��$X  H�D$�    �L$�L$D��1���@  1�H��$�   H�    H�$H��$P  H�\$H��$X  H�\$H��$�   H�\$�    �L$D�\$ �� ��   H��$�   H��$�   H��$�   H��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I������q���  1�H��$p  H��$x  H��$�  H��$�  H�    H�$H��$P  H�\$H��$X  H�\$H��$p  H�\$�    �\$ �� ��  H��$�   H��$�   H�    1�H9��T  H��$�   H��$p  H��$x  1�H��$�  H��$�  H��$   H��$  H�D$X    1�H��$�  H��$�  H��$�  H��$�  H��$0  H��$�  H��$8  H��$�  H�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�\$(H��$�  H�H�M H�KH�MH��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$   H��$�  H��$  H��$�  H��$p  H��$�  H��$x  H��$�  H��$�  H��$�  H��$�  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$P  H�\$0H��$X  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$P  H��$  H��$X  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H�D$�z���H�    H��$�  HǄ$�     H�    H�$H��$�  H�\$H�D$    �    H�\$H�H�$H�KH�L$�    =�Tu�H�D$P    H�    H�$H�T$H�L$H�\$PH�\$�    �\$ �� �a���H��$  H��$  H��$p  H�$H��$x  H�D$�    H��$p  H��$x  �L$���T��  �L$D��1���K  1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$p  H��$x  �L$D�\$ �� ��   H�\$PH�$�    H�\$H��$�   H��$�   H��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I������T�����H�D$H    H�    H�$H�l$H�T$H�\$HH�\$�    �\$ �� �q���H�\$PH�\$`H�\$HH�\$XH�    H�$H�    H�\$H�    H�\$H�\$`H�\$H�D$     �    H�\$(H��$p  H�\$0H��$x  H�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�L$(H�D$0H��$p  H��$  H��$x  H��$   H��$(  H��$0  H���  ÉL$D����>�K  1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$p  H��$x  �L$D�\$ �� ��   H�\$PH�$�    H�\$H��$�   H��$�   H��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I�����@��q�K  1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$p  H��$x  �L$D�\$ �� ��   H�\$PH�$�    H�\$H��$  H��$�   H��$   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$  H��$   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I������q�������1�H��$P  H��$X  H��$`  H��$h  H�    H�$H�l$H�T$H��$P  H�\$�    �\$ �� �v���H�\$PH�\$`H�    H�$H�    H�\$H�    H�\$H�\$`H�\$H�D$     �    H�L$(H�D$0H��$P  H��$X  1�H��$�  H��$�  H��$�  H��$�  H�D$`    1�H��$�  H��$�  H��$�  H��$�  H��$@  H��$�  H��$H  H��$�  H�    H�$H�    H�\$H�    H�\$H�\$`H�\$H�D$     �    H�\$(H��$�  H�H�M H�KH�MH��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$P  H��$�  H��$X  H��$�  H��$`  H��$�  H��$h  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$P  H�\$0H��$X  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$P  H��$  H��$X  H��$   H��$(  H��$0  H���  ÉD$D=��
&uyH�    H�$H�T$H�L$H�D$    �    H��$p  H��$x  �D$D�\$ �� t8H��$  H��$   H��$  H��$(  H��$  H��$0  H���  �=��>�L���1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    �\$ �� ����H��$  H��$  H��$P  H�$H��$X  H�D$�    �L$�L$D��1���N  1�H��$�   H�    H�$H��$P  H�\$H��$X  H�\$H��$�   H�\$�    �L$D�\$ �� ��   H��$�   H�$�    H�\$H��$�   H��$�   H��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I�������>�7  1�H�\$xH�    H�$H��$P  H�\$H��$X  H�\$H�\$xH�\$�    �L$D�\$ �� ��   H��$�   H��$�   H�\$xH��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I������q���.���1�H��$0  H��$8  H��$@  H��$H  H�    H�$H��$P  H�\$H��$X  H�\$H��$0  H�\$�    �\$ �� �����H��$�   H��$�   H�    1�H9��T  H��$�   H��$P  H��$X  1�H��$�  H��$�  H��$�  H��$�  H�D$X    1�H��$�  H��$�  H��$�  H��$�  H��$  H��$�  H��$  H��$�  H�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�\$(H��$�  H�H�M H�KH�MH��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$0  H��$�  H��$8  H��$�  H��$@  H��$�  H��$H  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$p  H�\$0H��$x  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$p  H��$  H��$x  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H�D$�z���=@��q��  �D$D=�|~?�  1�H�    H�$H�T$H�L$H�\$DH�\$�    H��$p  H��$x  �D$D�\$ �� ��   H�    H�$H�    H�\$H�    H�\$H�\$DH�\$H�D$     �    H�\$(H��$`  H�\$0H��$h  H�    H�$H�    H�\$H�    H�\$H�\$DH�\$H�D$     �    H�L$(H�D$0H��$`  H��$  H��$h  H��$   H��$(  H��$0  H���  �=@��q�����1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    �\$ �� �����H��$  H��$  H��$p  H�$H��$x  H�D$�    H��$p  H��$x  �L$����>��  �L$D��1���N  1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$p  H��$x  �L$D�\$ �� ��   H��$�   H�$�    H�\$H��$�   H��$�   H��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I�������>�����1�H�\$pH�    H�$H�l$H�T$H�\$pH�\$�    �\$ �� �����H��$�   H�$�    H�\$H��$�   H�\$pH��$�   H�5    H��$�   1�H9�t}H�    1�H9�t8H��$�   H��$�   H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I����L$D��@��q�@  1�H��$�   H�    H�$H�l$H�T$H��$�   H�\$�    H��$p  H��$x  �L$D�\$ �� ��   H��$�   H��$   H��$�   H��$  H�5    H��$�   1�H9�t}H�    1�H9�t8H��$   H��$  H��$  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H��$�   H�D$�H�    H�$H�    H�\$H�    H�\$�    H�t$H��$�   �I������q���\���1�H��$  H��$  H��$   H��$(  H�    H�$H�l$H�T$H��$  H�\$�    �\$ �� ����H��$�   H��$   H�    1�H9��T  H��$   H��$P  H��$X  1�H��$�  H��$�  H��$�  H��$�  H�D$`    1�H��$�  H��$�  H��$�  H��$�  H��$   H��$�  H��$(  H��$�  H�    H�$H�    H�\$H�    H�\$H�\$`H�\$H�D$     �    H�\$(H��$�  H�H�M H�KH�MH��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$  H��$�  H��$  H��$�  H��$   H��$�  H��$(  H��$�  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�\$(H��$p  H�\$0H��$x  H�    H�$H�    H�\$H�    H�\$H��$�  H�\$H�D$     �    H�L$(H�D$0H��$p  H��$  H��$x  H��$   H��$(  H��$0  H���  �H�    H�$H�    H�\$H�    H�\$�    H�D$�z����D$D=�n�uEH�    H�$H�T$H�L$H�D$    �    H��$p  H��$x  �D$D�\$ �� �~���=�q������H�    H�$H�T$H�L$H�D$    �    H��$p  H��$x  �\$ �� �2��������    �>������������������
      \�  runtime.duffzero   p�  runtime.duffzero   �  "".ord   �  "".ord   �  "".match   �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  $runtime.ifacethash   �   type."".floatVal   �	  $runtime.assertI2T2   �
  8go.itab."".floatVal."".Value   �
  8go.itab."".floatVal."".Value   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  $type."".complexVal   �  $runtime.assertI2T2   �  8go.itab."".floatVal."".Value   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �  $type."".complexVal   �  type."".Value   �  <go.itab."".complexVal."".Value   �  runtime.convT2I   �   type."".floatVal   �  type."".Value   �  8go.itab."".floatVal."".Value   �   runtime.typ2Itab   �  .go.string."unreachable"   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �   type."".int64Val   �  $runtime.assertI2T2   �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �  "".i64tof   �  8go.itab."".floatVal."".Value   �   8go.itab."".floatVal."".Value   �!   type."".floatVal   �!  type."".Value   �!  8go.itab."".floatVal."".Value   �!   runtime.typ2Itab   �"   type."".floatVal   �"  type."".Value   �"  8go.itab."".floatVal."".Value   �"   runtime.typ2Itab   �#   type."".int64Val   �#  $runtime.assertI2T2   �$   type."".int64Val   �$  type."".Value   �$  8go.itab."".int64Val."".Value   �%  runtime.convT2I   �%   type."".int64Val   �%  type."".Value   �&  8go.itab."".int64Val."".Value   �&  runtime.convT2I   �(  type."".ratVal   �(  $runtime.assertI2T2   �)  "".i64tor   �)  4go.itab."".ratVal."".Value   �*  4go.itab."".ratVal."".Value   �+  type."".ratVal   �+  type."".Value   �+  4go.itab."".ratVal."".Value   �+   runtime.typ2Itab   �,  type."".ratVal   �,  type."".Value   �,  4go.itab."".ratVal."".Value   �,   runtime.typ2Itab   �-  type."".intVal   �-  $runtime.assertI2T2   �.  "".i64toi   �/  4go.itab."".intVal."".Value   �/  4go.itab."".intVal."".Value   �0  type."".intVal   �0  type."".Value   �1  4go.itab."".intVal."".Value   �1   runtime.typ2Itab   �1  type."".intVal   �1  type."".Value   �1  4go.itab."".intVal."".Value   �2   runtime.typ2Itab   �3  $type."".complexVal   �3  $runtime.assertI2T2   �4   type."".int64Val   �4  type."".Value   �4  8go.itab."".int64Val."".Value   �4  runtime.convT2I   �7   type."".int64Val   �7  type."".Value   �7  8go.itab."".int64Val."".Value   �8  runtime.convT2I   �;  $type."".complexVal   �;  type."".Value   �;  <go.itab."".complexVal."".Value   �;  runtime.convT2I   �<  $type."".complexVal   �<  type."".Value   �<  <go.itab."".complexVal."".Value   �=  runtime.convT2I   �>  type."".boolVal   �?  $runtime.assertI2T2   �@  type."".ratVal   �A  $runtime.assertI2T2   �B  $runtime.ifacethash   �B   type."".floatVal   �C  $runtime.assertI2T2   �D  "".rtof   �D  8go.itab."".floatVal."".Value   �E  8go.itab."".floatVal."".Value   �F   type."".floatVal   �F  type."".Value   �F  8go.itab."".floatVal."".Value   �F   runtime.typ2Itab   �G   type."".floatVal   �G  type."".Value   �G  8go.itab."".floatVal."".Value   �G   runtime.typ2Itab   �H  type."".ratVal   �H  $runtime.assertI2T2   �I  4go.itab."".ratVal."".Value   �J  4go.itab."".ratVal."".Value   �K  type."".ratVal   �K  type."".Value   �K  4go.itab."".ratVal."".Value   �K   runtime.typ2Itab   �L  type."".ratVal   �L  type."".Value   �L  4go.itab."".ratVal."".Value   �L   runtime.typ2Itab   �M  $type."".complexVal   �N  $runtime.assertI2T2   �O  4go.itab."".ratVal."".Value   �Q   type."".int64Val   �Q  type."".Value   �Q  8go.itab."".int64Val."".Value   �R  runtime.convT2I   �U  $type."".complexVal   �U  type."".Value   �U  <go.itab."".complexVal."".Value   �V  runtime.convT2I   �V  $type."".complexVal   �V  type."".Value   �V  <go.itab."".complexVal."".Value   �W  runtime.convT2I   �X  type."".ratVal   �X  type."".Value   �X  4go.itab."".ratVal."".Value   �Y   runtime.typ2Itab   �Y  $type."".unknownVal   �Z  $runtime.assertI2T2   �Z  $type."".unknownVal   �[  type."".Value   �[  <go.itab."".unknownVal."".Value   �[  runtime.convT2I   �\  $type."".unknownVal   �\  type."".Value   �\  <go.itab."".unknownVal."".Value   �]  runtime.convT2I   �^  type."".intVal   �_  $runtime.assertI2T2   �_  $runtime.ifacethash   �`   type."".floatVal   �a  $runtime.assertI2T2   �b  "".itof   �b  8go.itab."".floatVal."".Value   �c  8go.itab."".floatVal."".Value   �d   type."".floatVal   �d  type."".Value   �d  8go.itab."".floatVal."".Value   �d   runtime.typ2Itab   �e   type."".floatVal   �e  type."".Value   �e  8go.itab."".floatVal."".Value   �e   runtime.typ2Itab   �f  type."".ratVal   �f  $runtime.assertI2T2   �g  "".itor   �g  4go.itab."".ratVal."".Value   �h  4go.itab."".ratVal."".Value   �i  type."".ratVal   �i  type."".Value   �i  4go.itab."".ratVal."".Value   �i   runtime.typ2Itab   �j  type."".ratVal   �j  type."".Value   �j  4go.itab."".ratVal."".Value   �j   runtime.typ2Itab   �k  type."".intVal   �k  $runtime.assertI2T2   �m  4go.itab."".intVal."".Value   �m  4go.itab."".intVal."".Value   �n  type."".intVal   �n  type."".Value   �n  4go.itab."".intVal."".Value   �n   runtime.typ2Itab   �o  type."".intVal   �o  type."".Value   �o  4go.itab."".intVal."".Value   �o   runtime.typ2Itab   �p  $type."".complexVal   �q  $runtime.assertI2T2   �r  4go.itab."".intVal."".Value   �t   type."".int64Val   �t  type."".Value   �t  8go.itab."".int64Val."".Value   �u  runtime.convT2I   �x  $type."".complexVal   �x  type."".Value   �x  <go.itab."".complexVal."".Value   �y  runtime.convT2I   �y  $type."".complexVal   �y  type."".Value   �y  <go.itab."".complexVal."".Value   �z  runtime.convT2I   �{  type."".intVal   �{  type."".Value   �{  4go.itab."".intVal."".Value   �|   runtime.typ2Itab   �|  "type."".stringVal   �}  $runtime.assertI2T2   �}  $type."".complexVal   �~  $runtime.assertI2T2   �~  0runtime.morestack_noctxt   ��  �"".autotmp_0604  type."".Value "".autotmp_0603  type."".Value "".autotmp_0602  $type."".complexVal "".autotmp_0601  type.*uint8 "".autotmp_0600  type."".Value "".autotmp_0599  type."".Value "".autotmp_0598  type."".Value "".autotmp_0597  type.*uint8 "".autotmp_0596  type.*uint8 "".autotmp_0595  type.uint32 "".autotmp_0594  type.bool "".autotmp_0593  type."".Value "".autotmp_0592  type."".Value "".autotmp_0591  type."".Value "".autotmp_0590  $type."".complexVal "".autotmp_0589  type.*uint8 "".autotmp_0588  type."".Value "".autotmp_0587  type."".Value "".autotmp_0586  type."".Value "".autotmp_0585  type.*uint8 "".autotmp_0584  type.*uint8 "".autotmp_0583  type."".Value "".autotmp_0582  type."".Value "".autotmp_0581  type.*uint8 "".autotmp_0580  type.*uint8 "".autotmp_0579  type.uint32 "".autotmp_0578  type.bool "".autotmp_0577  type."".Value "".autotmp_0576  type."".Value "".autotmp_0575  type."".Value "".autotmp_0574  $type."".complexVal "".autotmp_0573  type.*uint8 "".autotmp_0572  type."".Value "".autotmp_0571  type."".Value "".autotmp_0570  type."".Value "".autotmp_0569  type.*uint8 "".autotmp_0568  type.*uint8 "".autotmp_0567  type."".Value "".autotmp_0566  type."".Value "".autotmp_0565  type.*uint8 "".autotmp_0564  type.*uint8 "".autotmp_0563  type."".Value "".autotmp_0562  type."".Value "".autotmp_0561  type.*uint8 "".autotmp_0560  type.*uint8 "".autotmp_0559  type.uint32 "".autotmp_0558  type.bool "".autotmp_0557  type."".Value "".autotmp_0556  type."".Value "".autotmp_0555  type."".Value "".autotmp_0554 �$type."".complexVal "".autotmp_0553  type."".Value "".autotmp_0552  type."".Value "".autotmp_0551  type."".Value "".autotmp_0550  type.*uint8 "".autotmp_0549  type.*uint8 "".autotmp_0548  type."".Value "".autotmp_0547  type."".Value "".autotmp_0546  type.*uint8 "".autotmp_0545  type.*uint8 "".autotmp_0544  type."".Value "".autotmp_0543  type."".Value "".autotmp_0542 �type.*uint8 "".autotmp_0541 �type.*uint8 "".autotmp_0540  type."".Value "".autotmp_0539  type."".Value "".autotmp_0538  type.uint32 "".autotmp_0537  type.bool "".autotmp_0536  type."".Value "".autotmp_0535 �type."".Value "".autotmp_0534 �type."".Value "".autotmp_0533 �
type.uint32 "".autotmp_0531 �type."".Value "".autotmp_0530 �type.string "".autotmp_0529  $type."".complexVal "".autotmp_0528  $type."".complexVal "".autotmp_0527   type."".int64Val "".autotmp_0526   type."".floatVal "".autotmp_0525   type."".floatVal "".autotmp_0524   type."".floatVal "".autotmp_0523  $type."".complexVal "".autotmp_0522  $type."".complexVal "".autotmp_0521   type."".int64Val "".autotmp_0520  type."".ratVal "".autotmp_0519   type."".floatVal "".autotmp_0518   type."".floatVal "".autotmp_0517  type."".ratVal "".autotmp_0516  type."".ratVal "".autotmp_0515  $type."".complexVal "".autotmp_0514  $type."".complexVal "".autotmp_0513   type."".int64Val "".autotmp_0512  type."".intVal "".autotmp_0511   type."".floatVal "".autotmp_0510   type."".floatVal "".autotmp_0509  type."".ratVal "".autotmp_0508  type."".ratVal "".autotmp_0507  type."".intVal "".autotmp_0506  type."".intVal "".autotmp_0505 $type."".complexVal "".autotmp_0504 ?$type."".complexVal "".autotmp_0503   type."".int64Val "".autotmp_0502   type."".int64Val "".autotmp_0501 � type."".floatVal "".autotmp_0500 � type."".floatVal "".autotmp_0499 �type."".ratVal "".autotmp_0498 �type."".ratVal "".autotmp_0497 �type."".intVal "".autotmp_0496 �type."".intVal "".autotmp_0495 �
 type."".int64Val "".autotmp_0494 �
 type."".int64Val "".autotmp_0493 �
$type."".unknownVal "".autotmp_0492 �
$type."".unknownVal "".autotmp_0490 �
type.int "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".~r1 �$type."".complexVal "".x �type."".Value "".y �$type."".complexVal "".y �	 type."".floatVal "".x � type."".floatVal "".y �$type."".complexVal "".y �	 type."".floatVal "".y �	type."".ratVal "".x �type."".ratVal "".y �$type."".complexVal "".y �	 type."".floatVal "".y �	type."".ratVal "".y �	type."".intVal "".x �type."".intVal "".y �$type."".complexVal "".y � type."".floatVal "".y �	type."".ratVal "".y �	type."".intVal "".y �
 type."".int64Val "".x �
 type."".int64Val "".x �
$type."".unknownVal "".~b3 `type."".Value "".~b2 @type."".Value "".y  type."".Value "".x  type."".Value �"������������������������������������������������������ �? ��de<(�V��s�]eB��G�c�_�c�#L
8	JD��Y�s�Ob�J,��E�c�c�;�fs � }���7w��XjKP'<��7K���7O0�7g��Xp�<x�7Y�7w��XjJ]U ~<��7I�"7S�"7g��Xj8#� Tgclocals·7f2bc03eae9ababa8d2e476fa773c6e9 Tgclocals·6964cae77cc8ca448bf07954c3733ae6   @$GOROOT/src/go/constant/value.go�"".BinaryOp  �j  �jdH�%    H��$0���H;A��  H��P  W��$�  �$�  �$  �$�   �$�   1�H��$�  H��$�  H��$X  H�$H��$`  H�\$H��$p  H�\$H��$x  H�\$�    H�L$ H�D$(H�\$0H��$p  H�\$8H��$x  H��$X  H��$`  H��$  H�$H��$   H�D$�    H��$  H��$   �D$=��>��  =�T��  �D$D=1���  1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    H��$  H��$   �D$D�\$ �� ��  H��$�   H��$�   1�H��$�   H�    H�$H��$p  H�\$H��$x  H�\$H��$�   H�\$�    H��$�   H��$�   �    H��$�   H��$�   H�,$H��$h  H����  H��uNH��$�   H�,$H�T$H�L$�    H��$�   H�$�    H�L$H�D$H��$�  H��$�  H��P  �H��uH��$�   H�,$H�T$H�L$�    �H��$h  H�\$X1�H��$   H��$(  H��$0  H��$8  H��$@  H��$H  H��$   H�� �
  HǄ$�     HǄ$�     H��$�  H��$X  H�$H��$`  H�\$�    H�L$H�D$H��$�  H��$  H�H��$  �=     ��  H�CH�    H�$H�\$XH�\$H�D$    �    H�L$H�D$ H��$�  H��H��$  H�H��$  �=     �  H�CH��$p  H�$H��$x  H�\$�    H�L$H�D$H��$�  H�� H��$  H�H��$  �=     ��   H�CH�    H�$H�D$!   H��$�  H�\$H��$�  H�\$H��$�  H�\$ �    H�\$(H��$(  H�\$0H��$0  H�    H�$H��$(  H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M���L�CL�$H�D$�    �����L�CL�$H�D$�    �j���������H��u H��$�   H�,$H�T$H�L$�    �"���H���n���H��$�   H�,$H�T$H�L$�    �����=�T�C���H�D$H    H�    H�$H�T$H�L$H�\$HH�\$�    �\$ �� ����H�\$HH�\$hH�D$`    H�    H�$H��$p  H�\$H��$x  H�\$H�\$`H�\$�    H�L$hH�T$`H�T$PH��$h  H���}  H���  H���6  H�$�    �\$�� ��   H�\$PH�$�    �\$�� toH�L$hH�l$PH�H�L$`H�    H�$H�    H�\$H�    H�\$H�\$`H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H��P  �H�    H�$�    H�\$H�\$pH�\$hH�$�    H�\$H��$�   H�\$PH�$�    H�D$H�\$pH�$H��$�   H�\$H�D$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H��P  �H���L���H�$�    �\$�� t*H�\$PH�$�    �\$�� tH�L$hH�l$PH)�����H�    H�$�    H�\$H�\$xH�\$hH�$�    H�\$H��$�   H�\$PH�$�    H�D$H�\$xH�$H��$�   H�\$H�D$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H��P  �H����   H�$�    �\$�� t+H�\$PH�$�    �\$�� tH�L$hH�l$PH�������H�    H�$�    H�\$H��$�   H�\$hH�$�    H�\$H��$�   H�\$PH�$�    H�D$H��$�   H�$H��$�   H�\$H�D$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H��P  �H��u>H�$H�T$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H��P  �H���C���H��H��H���tH�H��H�������1������H�� H��uH!�����H������H	�����H��uH1�����H��uH��H���H!�H������H�������H��H��H���tH�H��H���d���H��H���Y����D$D=��
&�  �D$B H�    H�$H�T$H�L$H�\$BH�\$�    H��$  H��$   �D$D�\$ �� �4  �D$C H�    H�$H��$p  H�\$H��$x  H�\$H�\$CH�\$�    �\$CH��$h  H��"uo�|$B ta�\$CH�    H�$H�    H�\$H�    H�\$H�\$CH�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H��P  ��D$C �H��#������|$B ua�\$CH�    H�$H�    H�\$H�    H�\$H�\$CH�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H��P  ��D$C�=��>����1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    �\$ �� �����H��$�   H��$   1�H��$�   H�    H�$H��$p  H�\$H��$x  H�\$H��$�   H�\$�    H��$�   H��$�   H�    H�$�    H��$   H��$�   H�l$H��$h  H��{H��uNH��$�   H�,$H�T$H�L$�    H��$�   H�$�    H�L$H�D$H��$�  H��$�  H��P  �H�������H��$�   H�,$H�T$H�L$�    �H��uH��$�   H�,$H�T$H�L$�    �H�������H��$�   H�,$H�T$H�L$�    �Y���=@��q��  �D$D=�|~?��   1�H�    H�$H�T$H�L$H�\$BH�\$�    H��$  H��$   �D$D�\$ �� t]H�    H�$H�    H�\$H�    H�\$H�\$BH�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H��P  �=@��q�����1�H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    �\$ �� �p���H��$�   H��$�   1�H��$�   H�    H�$H��$p  H�\$H��$x  H�\$H��$�   H�\$�    H��$�   H��$�   H�    H�$�    H��$�   H��$�   H�l$H��$h  H���<  H��{H��uNH��$�   H�,$H�T$H�L$�    H��$�   H�$�    H�L$H�D$H��$�  H��$�  H��P  �H���t���H��$�   H�,$H�T$H�L$�    �H��uH��$�   H�,$H�T$H�L$�    �H��uhH�    H�$�    H�\$H�$H��$�   H�\$H��$�   H�\$�    H�\$H�$�    H�L$H�D$H��$�  H��$�  H��P  �H�������H��$�   H�,$H�T$H�L$�    �����H��PH��u H��$�   H�,$H�T$H�L$�    ����H���f���H��$�   H�,$H�T$H�L$�    ����H��u H��$�   H�,$H�T$H�L$�    �o���H��u H��$�   H�,$H�T$H�L$�    �I���H�������H��$�   H�,$H�T$H�L$�    �����D$D=�n��q  1�H��$  H��$   H�    H�$H�T$H�L$H��$  H�\$�    H��$  H��$   �D$D�\$ �� �  H��$h  H���T���1�H��$H  H��$P  H�    H�$H��$p  H�\$H��$x  H�\$H��$H  H�\$�    H�$    H��$  H�\$H��$   H�\$H��$H  H�\$H��$P  H�\$ �    H�\$(H��$8  H�\$0H��$@  H�    H�$H�    H�\$H�    H�\$H��$8  H�\$H�D$     �    H�\$(H��$�  H�\$0H��$�  H��P  �=�q���E���1�H��$�  H��$�  H��$�  H��$�  H�    H�$H�T$H�L$H��$�  H�\$�    �\$ �� �����1�H��$   H��$  H��$  H��$  H�    H�$H��$p  H�\$H��$x  H�\$H��$   H�\$�    L��$   L��$  H��$  H��$  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$�  H��$   H��$�  H��$�  L��$�  L��$�  L��$�  L��$�  H��$  H��$�  H��$   H��$�  1�H��$H  H��$P  1�H��$h  H��$p  H��$h  H����  H���h  H�4$H�l$L�L$L�D$�    H�\$ H��$H  H�\$(H��$P  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�L$ H�D$(H��$H  H��$P  H��$h  H��$p  1�H��$  H��$  1�H��$   H��$  H��$  H��$  H��$8  H��$   H��$@  H��$  H��$X  H��$  H��$`  H��$  H�    H�$H�    H�\$H�    H�\$H��$   H�\$H�D$     �    H�L$(H�D$0H��$�  H��$�  H��P  �H���3���H�4$H�l$L�L$L�D$�    H�\$ H��$H  H�\$(H��$P  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�L$ H�D$(����H����  H�4$H�l$L�L$L�D$�    H�\$ H��$x  H�\$(H��$�  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$�  H�\$(H��$�  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$�  H�\$(H��$�  H��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$X  H�\$(H��$`  H��$x  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$H  H�\$(H��$P  H��$�  H�$H��$�  H�\$H��$X  H�\$H��$`  H�\$�    H�L$ H�D$(����H�������H�4$H�l$L�L$L�D$�    H�\$ H��$�  H�\$(H��$�  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$�  H�\$(H��$�  H��$�  H�$H��$   H�\$H��$�  H�\$H��$�  H�\$�    H�\$ H��$�  H�\$(H��$�  H��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H��$�  H��$�  H�\$ H��$h  H�\$(H��$p  H�$H�D$H�L$H�D$�    H��$�  H��$�  H�\$ H��$�  H�\$(H��$�  H�$H�D$H�L$H�D$�    H�L$ H�D$(H��$�  H�$H��$�  H�\$H��$x  H�L$H��$�  H�D$�    H�\$ H��$(  H�\$(H��$0  H��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�L$ H�D$(H��$H  H�$H��$P  H�D$H��$(  H�\$H��$0  H�\$�    H�\$ H��$H  H�\$(H��$P  H��$�  H�$H��$�  H�\$H��$h  H�\$H��$p  H�\$�    H�L$ H�D$(H��$h  H�$H��$p  H�D$H��$(  H�\$H��$0  H�\$�    H�L$ H�D$(�����    �X����������̬
      �  "".match   �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".floatVal   �  "runtime.assertI2T   �  "".newFloat   �  *math/big.(*Float).Add   �  "".makeFloat   �	  *math/big.(*Float).Sub   �  runtime.convI2E   � (runtime.writeBarrier   �  &type.go/token.Token   �  runtime.convT2E   � (runtime.writeBarrier   �  runtime.convI2E   � (runtime.writeBarrier   �  Zgo.string."invalid binary operation %v %s %v"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  *math/big.(*Float).Mul   �  *math/big.(*Float).Quo   �   type."".int64Val   �  $runtime.assertI2T2   �   type."".int64Val   �  "runtime.assertI2T   �  "".is63bit   �  "".is63bit   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "type.math/big.Int   �  "runtime.newobject   �  math/big.NewInt   �  math/big.NewInt   �  &math/big.(*Int).Add   �  "".makeInt   �  "".is63bit   �  "".is63bit   �  "type.math/big.Int   �  "runtime.newobject   �  math/big.NewInt   �  math/big.NewInt   �  &math/big.(*Int).Sub   �  "".makeInt   �   "".is32bit   �   "".is32bit   �!  "type.math/big.Int   �!  "runtime.newobject   �!  math/big.NewInt   �"  math/big.NewInt   �"  &math/big.(*Int).Mul   �#  "".makeInt   �#  math/big.NewRat   �$  "".makeRat   �'  type."".boolVal   �(  $runtime.assertI2T2   �(  type."".boolVal   �)  "runtime.assertI2T   �*  type."".boolVal   �*  type."".Value   �*  6go.itab."".boolVal."".Value   �*  runtime.convT2I   �+  type."".boolVal   �,  type."".Value   �,  6go.itab."".boolVal."".Value   �,  runtime.convT2I   �-  type."".ratVal   �.  $runtime.assertI2T2   �/  type."".ratVal   �/  "runtime.assertI2T   �0  "type.math/big.Rat   �0  "runtime.newobject   �1  &math/big.(*Rat).Add   �1  "".makeRat   �2  &math/big.(*Rat).Sub   �3  &math/big.(*Rat).Mul   �3  &math/big.(*Rat).Quo   �4  $type."".unknownVal   �4  $runtime.assertI2T2   �5  $type."".unknownVal   �5  type."".Value   �5  <go.itab."".unknownVal."".Value   �6  runtime.convT2I   �7  type."".intVal   �7  $runtime.assertI2T2   �8  type."".intVal   �9  "runtime.assertI2T   �9  "type.math/big.Int   �9  "runtime.newobject   �;  &math/big.(*Int).Add   �;  "".makeInt   �<  &math/big.(*Int).Sub   �<  &math/big.(*Int).Mul   �=  "type.math/big.Rat   �=  "runtime.newobject   �=  .math/big.(*Rat).SetFrac   �>  "".makeRat   �?  &math/big.(*Int).Rem   �?  &math/big.(*Int).And   �@  $math/big.(*Int).Or   �A  &math/big.(*Int).Xor   �A  ,math/big.(*Int).AndNot   �B  &math/big.(*Int).Quo   �C  "type."".stringVal   �C  $runtime.assertI2T2   �D  "type."".stringVal   �E  "runtime.assertI2T   �F  *runtime.concatstring2   �G  "type."".stringVal   �G  type."".Value   �G  :go.itab."".stringVal."".Value   �H  runtime.convT2I   �I  $type."".complexVal   �I  $runtime.assertI2T2   �J  $type."".complexVal   �K  "runtime.assertI2T   �O  "".add   �P  "".add   �S  $type."".complexVal   �S  type."".Value   �S  <go.itab."".complexVal."".Value   �T  runtime.convT2I   �U  "".sub   �V  "".sub   �W  "".mul   �X  "".mul   �Z  "".mul   �[  "".mul   �\  "".sub   �]  "".add   �^  "".mul   �_  "".mul   �a  "".mul   �b  "".mul   �c  "".mul   �d  "".mul   �e  "".add   �f  "".add   �g  "".quo   �i  "".sub   �j  "".quo   �j  0runtime.morestack_noctxt   p�  �"".autotmp_0690  "type.interface {} "".autotmp_0689  "type.interface {} "".autotmp_0688 �"type.interface {} "".autotmp_0687 _(type.[3]interface {} "".autotmp_0684 �&type.[]interface {} "".autotmp_0683  type."".Value "".autotmp_0682  &type.go/token.Token "".autotmp_0681  type."".Value "".autotmp_0680  type."".Value "".autotmp_0679  &type.go/token.Token "".autotmp_0678  &type.go/token.Token "".autotmp_0677  &type.go/token.Token "".autotmp_0676  &type.go/token.Token "".autotmp_0674 �type.uint32 "".autotmp_0672 �type."".Value "".autotmp_0671 �type.string "".autotmp_0670 �&type.go/token.Token "".autotmp_0669 �"type."".stringVal "".autotmp_0668 �"type."".stringVal "".autotmp_0667  $type."".complexVal "".autotmp_0666 �$type."".complexVal "".autotmp_0665  type."".Value "".autotmp_0664 �	 type."".floatVal "".autotmp_0663  type."".Value "".autotmp_0662  $type.*math/big.Rat "".autotmp_0661 �	type."".ratVal "".autotmp_0660  type."".Value "".autotmp_0659  type."".Value "".autotmp_0658  $type.*math/big.Rat "".autotmp_0657  $type.*math/big.Rat "".autotmp_0656  $type.*math/big.Int "".autotmp_0655 �	type."".intVal "".autotmp_0654   type."".int64Val "".autotmp_0653  type."".Value "".autotmp_0651  type."".Value "".autotmp_0650  $type.*math/big.Int "".autotmp_0649  $type.*math/big.Int "".autotmp_0648  $type.*math/big.Int "".autotmp_0647  $type.*math/big.Int "".autotmp_0646  type.bool "".autotmp_0645  type.bool "".autotmp_0644  type."".Value "".autotmp_0643  $type.*math/big.Int "".autotmp_0642  $type.*math/big.Int "".autotmp_0641  $type.*math/big.Int "".autotmp_0640  $type.*math/big.Int "".autotmp_0639  type.bool "".autotmp_0638  type.bool "".autotmp_0637  type."".Value "".autotmp_0636  $type.*math/big.Int "".autotmp_0634  $type.*math/big.Int "".autotmp_0633 �	$type.*math/big.Int "".autotmp_0631  type.bool "".autotmp_0630 � type."".int64Val "".autotmp_0629  type."".boolVal "".autotmp_0628  type."".boolVal "".autotmp_0627 �type."".boolVal "".autotmp_0626 �$type."".unknownVal "".~r2 �	type."".Value 
"".im �type."".Value 
"".re �type."".Value "".~r0 �$type.*math/big.Int "".~r0 �$type.*math/big.Int "".~r0 �$type.*math/big.Int "".x �"type."".stringVal "".s �type."".Value 
"".dd �type."".Value 
"".cc �type."".Value 
"".ad �type."".Value 
"".bc �type."".Value 
"".bd �type."".Value 
"".ac �type."".Value 
"".ad �type."".Value 
"".bc �type."".Value 
"".bd �type."".Value 
"".ac �type."".Value 
"".im �type."".Value 
"".re �type."".Value "".d �type."".Value "".c �type."".Value "".b �type."".Value "".a �type."".Value "".y �$type."".complexVal "".x �$type."".complexVal "".c �
(type.*math/big.Float "".b �
(type.*math/big.Float "".a �	(type.*math/big.Float "".x �
 type."".floatVal "".c �
$type.*math/big.Rat "".b �
$type.*math/big.Rat "".a �	$type.*math/big.Rat "".x �
type."".ratVal "".c �
$type.*math/big.Int "".b �
$type.*math/big.Int "".a �	$type.*math/big.Int "".x �type."".intVal "".b �type.int64 "".a �type.int64 "".x � type."".int64Val "".x �type."".boolVal "".x �$type."".unknownVal "".~r3 Ptype."".Value "".y 0type."".Value 
"".op  &type.go/token.Token "".x  type."".Value �"����������������C�����x���������������������
� �5 ��_\��Q3b�o	
�F
L
/8b;�
+.1�
+$'�>
A,
	
cZ
>o
oJ�Q%3
	
�^]JjQ%,3)
(%$!h
/
	
�j���b�y@P$
2B:�7
2B2/
2RRRRB"
2RRbB"RBRBB� � �R�GC�>�@.[=g�
%�%�(�[� DG�Y� NG ;(U �} �v#g&�R�DR1RRRRR	1R
RRBBBR�B& Tgclocals·4dd66991891153e33d6808f41376a850 Tgclocals·bbced691e09928f29a52c25e48674f8c   @$GOROOT/src/go/constant/value.go�"".add  �  �dH�%    H;av^H��81�H�\$`H�\$hH�\$@H�$H�\$HH�\$H�D$   H�\$PH�\$H�\$XH�\$ �    H�L$(H�D$0H�L$`H�D$hH��8��    �������������
      �  "".BinaryOp   �  0runtime.morestack_noctxt   `p  "".~r2 @type."".Value "".y  type."".Value "".x  type."".Value pYo � 
�� 
 O1 Tgclocals·8ead428b4183a0f1b19d8f59d3dde163 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".sub  �  �dH�%    H;av^H��81�H�\$`H�\$hH�\$@H�$H�\$HH�\$H�D$   H�\$PH�\$H�\$XH�\$ �    H�L$(H�D$0H�L$`H�D$hH��8��    �������������
      �  "".BinaryOp   �  0runtime.morestack_noctxt   `p  "".~r2 @type."".Value "".y  type."".Value "".x  type."".Value pYo � 
�� 
 O1 Tgclocals·8ead428b4183a0f1b19d8f59d3dde163 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".mul  �  �dH�%    H;av^H��81�H�\$`H�\$hH�\$@H�$H�\$HH�\$H�D$   H�\$PH�\$H�\$XH�\$ �    H�L$(H�D$0H�L$`H�D$hH��8��    �������������
      �  "".BinaryOp   �  0runtime.morestack_noctxt   `p  "".~r2 @type."".Value "".y  type."".Value "".x  type."".Value pYo � 
�� 
 O1 Tgclocals·8ead428b4183a0f1b19d8f59d3dde163 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".quo  �  �dH�%    H;av^H��81�H�\$`H�\$hH�\$@H�$H�\$HH�\$H�D$   H�\$PH�\$H�\$XH�\$ �    H�L$(H�D$0H�L$`H�D$hH��8��    �������������
      �  "".BinaryOp   �  0runtime.morestack_noctxt   `p  "".~r2 @type."".Value "".y  type."".Value "".x  type."".Value pYo � 
�� 
 O1 Tgclocals·8ead428b4183a0f1b19d8f59d3dde163 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�"".Shift  �  �dH�%    H�D$�H;A��  H���   1�H�D$`1�H��$  H��$  H��$�   H��$�   H��$�   H�$H��$�   H�D$�    H��$  �l$�l$<���T�	  H�D$@    H�    H�$H��$�   H�\$H��$�   H�\$H�\$@H�\$�    �l$<H��$  �\$ �� ��  H�� ugH�\$@H�\$XH�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�\$(H��$  H�\$0H��$  H���   �H��$   H��u^H�\$@H�$�    H�D$H�$H�D$H��$  H�\$�    H�\$H�$�    H�L$H�D$H��$  H��$  H���   �H��uyH�l$@H��H��@seH��H�l$XH�    H�$H�    H�\$H�    H�\$H�\$XH�\$H�D$     �    H�\$(H��$  H�\$0H��$  H���   �H��?�H��$   H�\$PH�T$H1�H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   H�� ��  HǄ$�      HǄ$�      H��$�   H��$�   H�$H��$�   H�\$�    H�L$H�D$H��$�   H�L$pH�H�D$x�=     �|  H�CH�    H�$H�\$PH�\$H�D$    �    H�L$H�D$ H��$�   H��H�L$pH�H�D$x�=     �  H�CH�    H�$H�\$HH�\$H�D$    �    H�L$H�D$ H��$�   H�� H�L$pH�H�D$x�=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$�   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M���L�CL�$H�D$�    �����L�CL�$H�D$�    �q������������|~?��   1�H�    H�$H��$�   H�\$H��$�   H�\$H�\$<H�\$�    �l$<H��$  �\$ �� t]H�    H�$H�    H�\$H�    H�\$H�\$<H�\$H�D$     �    H�\$(H��$  H�\$0H��$  H���   Á�@��q�����1�H�\$`H�    H�$H��$�   H�\$H��$�   H�\$H�\$`H�\$�    H��$  �\$ �� �����H�� udH�\$`H�\$hH�    1�H9�tH�\$hH��$  H��$  H���   �H�    H�$H�    H�\$H�    H�\$�    H�D$�H�    H�$�    H��$  H�D$H��$   H��uHH�$H�\$`H�\$H�T$�    H�\$H�$�    H�L$H�D$H��$  H��$  H���   �H�������H�$H�\$`H�\$H�T$�    H�\$H�$�    H�L$H�D$H��$  H��$  H���   ��    �*�������������f
      �  $runtime.ifacethash   �   type."".int64Val   �  $runtime.assertI2T2   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  "".i64toi   �  &math/big.(*Int).Lsh   �  "".makeInt   �   type."".int64Val   �  type."".Value   �  8go.itab."".int64Val."".Value   �  runtime.convT2I   �  runtime.convI2E   � (runtime.writeBarrier   �  &type.go/token.Token   �  runtime.convT2E   � (runtime.writeBarrier   �  type.uint   �  runtime.convT2E   � (runtime.writeBarrier   �  Dgo.string."invalid shift %v %s %d"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $type."".unknownVal   �  $runtime.assertI2T2   �  $type."".unknownVal   �  type."".Value   �  <go.itab."".unknownVal."".Value   �  runtime.convT2I   �  type."".intVal   �  $runtime.assertI2T2   �  4go.itab."".intVal."".Value   �  type."".intVal   �  type."".Value   �  4go.itab."".intVal."".Value   �   runtime.typ2Itab   �  "type.math/big.Int   �  "runtime.newobject   �  &math/big.(*Int).Lsh   �  "".makeInt   �  &math/big.(*Int).Rsh   �  "".makeInt   �  0runtime.morestack_noctxt   `�  :"".autotmp_0722  "type.interface {} "".autotmp_0721  "type.interface {} "".autotmp_0720 �"type.interface {} "".autotmp_0719 _(type.[3]interface {} "".autotmp_0716 �&type.[]interface {} "".autotmp_0715  &type.go/token.Token "".autotmp_0712 �type.uint32 "".autotmp_0710 �type."".Value "".autotmp_0709 �type.string "".autotmp_0708 �type.uint "".autotmp_0707 �&type.go/token.Token "".autotmp_0706  type."".Value "".autotmp_0705  $type.*math/big.Int "".autotmp_0704  type."".Value "".autotmp_0703  $type.*math/big.Int "".autotmp_0702  $type.*math/big.Int "".autotmp_0701  type."".intVal "".autotmp_0700   type."".int64Val "".autotmp_0699  type."".Value "".autotmp_0697 �type."".intVal "".autotmp_0696 � type."".int64Val "".autotmp_0695 �$type."".unknownVal "".x �type."".intVal "".x � type."".int64Val "".x �$type."".unknownVal "".~r3 @type."".Value "".s 0type.uint 
"".op  &type.go/token.Token "".x  type."".Value b����k��x�����������Q� � d�8�
gKy �9X]]"dH
H3 8 a���@.|Q�� Tgclocals·0588ca1c52d0ec7f6ca12931a37dd289 Tgclocals·4b6ac10bfefaa8263abce44bdd57d854   @$GOROOT/src/go/constant/value.go�"".cmpZero  �  �dH�%    H;a��   H��8H�L$@H�D$HH��)��   H��'uH�� �D$PH��8�H��(uH�� �D$PH��8�H��)uH�� �D$PH��8�H�    H�\$(H�D$0   H�    H�$H�\$(H�\$H�D$    �    H�\$H�H�$H�KH�L$�    H��,uH�� �D$PH��8�H��-uH�� �D$PH��8�H��.�z���H�� �D$PH��8��    ����������������
      �  .go.string."unreachable"   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  0runtime.morestack_noctxt   0p  "".autotmp_0724 type.string "".~r2  type.bool 
"".op &type.go/token.Token "".x  type.int 6p'opopopgopopo � D�T
  �v Tgclocals·f56b2291fa344104975cb6587be42b9b Tgclocals·d8fdd2a55187867c76648dc792366181   @$GOROOT/src/go/constant/value.go�"".Compare  �4  �4dH�%    H��$����H;A�  H��  W��$(  �$8  �$�   D$`D$hH��$�  H�$H��$�  H�\$H��$�  H�\$H��$�  H�\$�    H�L$ H�D$(H�\$0H��$�  H�\$8H��$�  H��$�  H��$�  H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �D$=��>�M  =�T��  �D$D=1����   1�H�\$hH�    H�$H�T$H�L$H�\$hH�\$�    H��$�   H��$�   �D$D�\$ �� ��   1�H�\$xH�    H�$H��$�  H�\$H��$�  H�\$H�\$xH�\$�    H�\$hH�$H�\$xH�\$�    H�\$H�$H��$�  H�\$�    �\$��$�  H�Ę  �=�T��   H�D$H    H�    H�$H�T$H�L$H�\$HH�\$�    �\$ �� ��   H�D$X    H�    H�$H��$�  H�\$H��$�  H�\$H�\$XH�\$�    H�L$XH��$�  H��)��  H��'uH�\$HH9���$�  H�Ę  �H��(uH�\$HH9���$�  H�Ę  �H��)uH�\$HH9���$�  H�Ę  �H��$�  H�\$P1�H��$h  H��$p  H��$x  H��$�  H��$�  H��$�  H��$h  H�� �
  HǄ$�      HǄ$      H��$�   H��$�  H�$H��$�  H�\$�    H�L$H�D$H��$�   H��$�   H�H��$�   �=     ��  H�CH�    H�$H�\$PH�\$H�D$    �    H�L$H�D$ H��$�   H��H��$�   H�H��$�   �=     �  H�CH��$�  H�$H��$�  H�\$�    H�L$H�D$H��$�   H�� H��$�   H�H��$�   �=     ��   H�CH�    H�$H�D$   H��$�   H�\$H��$�   H�\$H��$   H�\$ �    H�\$(H��$�   H�\$0H��$�   H�    H�$H��$�   H�\$H�D$    �    H�\$H�H�$H�KH�L$�    L�CL�$H�D$�    �M���L�CL�$H�D$�    �����L�CL�$H�D$�    �j���������H��,uH�\$HH9���$�  H�Ę  �H��-uH�\$HH9���$�  H�Ę  �H��.�X���H�\$HH9���$�  H�Ę  ÉD$D=��
&��   �D$A H�    H�$H�T$H�L$H�\$AH�\$�    H��$�   H��$�   �D$D�\$ �� ��   �D$C H�    H�$H��$�  H�\$H��$�  H�\$H�\$CH�\$�    �\$CH��H��$�  H��'u�\$A8���$�  H�Ę  �H��,�v����\$A8���$�  H�Ę  �=��>�T���1�H�\$`H�    H�$H�T$H�L$H�\$`H�\$�    �\$ �� ����1�H��$�   H�    H�$H��$�  H�\$H��$�  H�\$H��$�   H�\$�    H�\$`H�$H��$�   H�\$�    H�\$H�$H��$�  H�\$�    �\$��$�  H�Ę  �=@��q�.  �D$D=�|~?uT1�H�    H�$H�T$H�L$H�\$AH�\$�    H��$�   H��$�   �D$D�\$ �� tƄ$�   H�Ę  �=@��q����1�H�\$pH�    H�$H�T$H�L$H�\$pH�\$�    �\$ �� �����1�H��$�   H�    H�$H��$�  H�\$H��$�  H�\$H��$�   H�\$�    H�\$pH�$H��$�   H�\$�    H�\$H�$H��$�  H�\$�    �\$��$�  H�Ę  ÉD$D=�n���  1�H��$�   H��$�   H�    H�$H�T$H�L$H��$�   H�\$�    H��$�   H��$�   �D$D�\$ �� �X  1�H��$�   H��$�   H�    H�$H��$�  H�\$H��$�  H�\$H��$�   H�\$�    H��$�   H��$�   H��$�   H��$�   H��$�  H��)��   H��'uSH��$�   H9�u<H��$�   H�$H��$�   H�\$H�T$H�D$�    �\$ ��$�  H�Ę  �Ƅ$�   ��H��(uAH��$�   H�,$H��$�   H�l$H�T$H�D$�    H�\$ H�� ��$�  H�Ę  �H��)�����H��$�   H�,$H��$�   H�l$H�T$H�D$�    H�\$ H�� ��$�  H�Ę  �H��,uZH��$�   H9�uCH��$�   H�$H��$�   H�\$H�T$H�D$�    �\$ H��H����$�  H�Ę  �Ƅ$�  ��H��-uAH��$�   H�,$H��$�   H�l$H�T$H�D$�    H�\$ H�� ��$�  H�Ę  �H��.�����H��$�   H�,$H��$�   H�l$H�T$H�D$�    H�\$ H�� ��$�  H�Ę  �=�q�������1�H��$(  H��$0  H��$8  H��$@  H�    H�$H�T$H�L$H��$(  H�\$�    �\$ �� �3���1�H��$H  H��$P  H��$X  H��$`  H�    H�$H��$�  H�\$H��$�  H�\$H��$H  H�\$�    H��$H  H��$  H��$P  H��$  H��$X  H��$  H��$`  H��$   H��$(  H�H�$H�KH�L$H�D$'   H��$  H�|$H�H�H�KH�O�    �\$(�\$BH��$8  H�H�$H�KH�L$H�D$'   H��$  H�|$H�H�H�KH�O�    �T$B�\$(H��$�  H��H��'u�� t��$�  H�Ę  �Ƅ$�   ��H��,������� tH����$�  H�Ę  �Ƅ$�  ���    ��������~
      �  "".match   �  $runtime.ifacethash   �   type."".floatVal   �  $runtime.assertI2T2   �   type."".floatVal   �  "runtime.assertI2T   �  *math/big.(*Float).Cmp   �  "".cmpZero   �   type."".int64Val   �  $runtime.assertI2T2   �   type."".int64Val   �	  "runtime.assertI2T   �  runtime.convI2E   � (runtime.writeBarrier   �  &type.go/token.Token   �  runtime.convT2E   � (runtime.writeBarrier   �  runtime.convI2E   � (runtime.writeBarrier   �  Ngo.string."invalid comparison %v %s %v"   �  fmt.Sprintf   �  type.string   �  runtime.convT2E   �  runtime.gopanic   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  type."".boolVal   �  $runtime.assertI2T2   �  type."".boolVal   �  "runtime.assertI2T   �  type."".ratVal   �  $runtime.assertI2T2   �  type."".ratVal   �  "runtime.assertI2T   �  &math/big.(*Rat).Cmp   �  "".cmpZero   �  $type."".unknownVal   �  $runtime.assertI2T2   �  type."".intVal   �  $runtime.assertI2T2   �  type."".intVal   �   "runtime.assertI2T   �!  &math/big.(*Int).Cmp   �!  "".cmpZero   �"  "type."".stringVal   �"  $runtime.assertI2T2   �#  "type."".stringVal   �$  "runtime.assertI2T   �&   runtime.eqstring   �'  "runtime.cmpstring   �(  "runtime.cmpstring   �)   runtime.eqstring   �+  "runtime.cmpstring   �,  "runtime.cmpstring   �-  $type."".complexVal   �.  $runtime.assertI2T2   �.  $type."".complexVal   �/  "runtime.assertI2T   �1  "".Compare   �2  "".Compare   �4  0runtime.morestack_noctxt   `�  N"".autotmp_0754  "type.interface {} "".autotmp_0753  "type.interface {} "".autotmp_0752 �"type.interface {} "".autotmp_0751 _(type.[3]interface {} "".autotmp_0748 �&type.[]interface {} "".autotmp_0747  &type.go/token.Token "".autotmp_0746  &type.go/token.Token "".autotmp_0745  &type.go/token.Token "".autotmp_0743 �type.uint32 "".autotmp_0741 �type."".Value "".autotmp_0740 �type.string "".autotmp_0739 �&type.go/token.Token "".autotmp_0738 �"type."".stringVal "".autotmp_0737 �$type."".complexVal "".autotmp_0736  type.bool "".autotmp_0735  type.int "".autotmp_0734 � type."".floatVal "".autotmp_0733  type.bool "".autotmp_0732  type.int "".autotmp_0731 �type."".ratVal "".autotmp_0730  type.bool "".autotmp_0728 �type."".intVal "".autotmp_0727 � type."".int64Val "".autotmp_0726 �type."".boolVal "".y �"type."".stringVal "".x �"type."".stringVal 
"".re �type.bool "".y �$type."".complexVal "".x �$type."".complexVal "".x � type."".floatVal "".x �type."".ratVal "".x �type."".intVal "".x � type."".int64Val "".x �type."".boolVal "".x �$type."".unknownVal "".~r3 Ptype.bool "".y 0type."".Value 
"".op  &type.go/token.Token "".x  type."".Value �"����������������!����� �����i��������P��J��U��P��J�����+��
� � ��G\�J�IFBV�c
5Z
A
DD�CZD>�=jfiSA
AZA
AbP�JK
"c h zR���@.�[��dO�km	��Jw Tgclocals·8348f4c3fb43d484332abd834bc6b74d Tgclocals·5ea1f2fbb7a4500b5337d2bd0531ab03   @$GOROOT/src/go/constant/value.go�"".init  �  �dH�%    H;a�	  H���    �� t�    ��uH����    �    �    �    �    �    �    H�       �H�$�    H�\$�=     ��   H�    H��������H�$�    H�\$�=     uCH�    �    H�$�=     uH�    �    H���H�-    H�,$H�\$�    ��H�-    H�,$H�\$�    �H�-    H�,$H�\$�    �k����    ���������������6
      4  "".initdone·   L  "".initdone·   j  "runtime.throwinit   z "".initdone·   �  fmt.init   �  go/token.init   �  math.init   �  math/big.init   �  strconv.init   �  math/big.NewInt   � (runtime.writeBarrier   �  "".minInt64   �  math/big.NewInt   � (runtime.writeBarrier   �  "".maxInt64   �  "".newFloat   � (runtime.writeBarrier   �  "".floatVal0   � "".initdone·   �  "".floatVal0   �  .runtime.writebarrierptr   �  "".maxInt64   �  .runtime.writebarrierptr   �  "".minInt64   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt           � H � @�[�,(6����67�  4� Tgclocals·33cdeccccebe80329f1fdbee7f5874cb Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�$"".(*boolVal).Kind  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  &go.string."boolVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this   type.*"".boolVal `_`	_ � � 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�("".(*boolVal).String  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$8�+1�1�@�� tH�    H��   H�L$@H�D$HH��0�H�    H��   ���    �7����������
      |  (go.string."constant"   �  &go.string."boolVal"   �  $go.string."String"   �  "runtime.panicwrap   �   go.string."true"   �  "go.string."false"   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this   type.*"".boolVal `�_`_ � � 
 yW Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�2"".(*boolVal).ExactString  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$8�+1�1�1�@�� tH�    H��   H�L$@H�D$HH��0�H�    H��   ���    �5��������
      |  (go.string."constant"   �  &go.string."boolVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �   go.string."true"   �  "go.string."false"   �  0runtime.morestack_noctxt   0`  "".autotmp_0762  type.string "".~r0 type.string ""..this   type.*"".boolVal `�_`_ � � 
 yW Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�:"".(*boolVal).implementsValue  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  &go.string."boolVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this   type.*"".boolVal `s_`	_ � 
� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�("".(*stringVal).Kind  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  *go.string."stringVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  $type.*"".stringVal `_`	_ � � 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�,"".(*stringVal).String  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�t$8H�H�$H�NH�L$�    H�L$H�D$H�L$@H�D$HH��0��    �9������������
      �  (go.string."constant"   �  *go.string."stringVal"   �  $go.string."String"   �  "runtime.panicwrap   �  &"".stringVal.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  $type.*"".stringVal `�_ � �  �M Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�6"".(*stringVal).ExactString  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�t$8H�H�$H�NH�L$�    H�L$H�D$H�L$@H�D$HH��0��    �9������������
      �  (go.string."constant"   �  *go.string."stringVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  0"".stringVal.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  $type.*"".stringVal `�_ � �  �M Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�>"".(*stringVal).implementsValue  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  *go.string."stringVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  $type.*"".stringVal `s_`	_ � � 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�&"".(*int64Val).Kind  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  (go.string."int64Val"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  "type.*"".int64Val `_`	_ � � 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�*"".(*int64Val).String  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$8H�+H�,$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  (go.string."int64Val"   �  $go.string."String"   �  "runtime.panicwrap   �  $"".int64Val.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  "type.*"".int64Val `�_ � �  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�4"".(*int64Val).ExactString  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$8H�+H�,$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  (go.string."int64Val"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  ."".int64Val.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  "type.*"".int64Val `�_ � �  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�<"".(*int64Val).implementsValue  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  (go.string."int64Val"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  "type.*"".int64Val `s_`	_ � � 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�""".(*intVal).Kind �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  $go.string."intVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  type.*"".intVal `_`	_ � � 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�&"".(*intVal).String �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  $go.string."intVal"   �  $go.string."String"   �  "runtime.panicwrap   �   "".intVal.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  type.*"".intVal `�_ � �  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�0"".(*intVal).ExactString �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  $go.string."intVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  *"".intVal.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  type.*"".intVal `�_ �  �  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�8"".(*intVal).implementsValue �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  $go.string."intVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  type.*"".intVal `s_`	_ � "� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�""".(*ratVal).Kind �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  $go.string."ratVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  type.*"".ratVal `_`	_ � $� 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�&"".(*ratVal).String �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  $go.string."ratVal"   �  $go.string."String"   �  "runtime.panicwrap   �   "".ratVal.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  type.*"".ratVal `�_ � &�  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�0"".(*ratVal).ExactString �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  $go.string."ratVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  *"".ratVal.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  type.*"".ratVal `�_ � (�  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�8"".(*ratVal).implementsValue �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  $go.string."ratVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  type.*"".ratVal `s_`	_ � *� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�&"".(*floatVal).Kind �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  (go.string."floatVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  "type.*"".floatVal `_`	_ � ,� 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�*"".(*floatVal).String �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  (go.string."floatVal"   �  $go.string."String"   �  "runtime.panicwrap   �  $"".floatVal.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  "type.*"".floatVal `�_ � .�  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�4"".(*floatVal).ExactString �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�t$8H�H�$�    H�L$H�D$H�L$@H�D$HH��0��    �B�����
      �  (go.string."constant"   �  (go.string."floatVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  ."".floatVal.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  "type.*"".floatVal `�_ � 0�  �= Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�<"".(*floatVal).implementsValue �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  (go.string."floatVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  "type.*"".floatVal `s_`	_ � 2� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�4type..hash.[1]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0774 type.int "".autotmp_0773 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[1]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�0type..eq.[1]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0778 ?"type.interface {} "".autotmp_0777 "type.interface {} "".autotmp_0776 _type.int "".autotmp_0775 Otype.int "".~r2  type.bool "".q *type.*[1]interface {} "".p  *type.*[1]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   @$GOROOT/src/go/constant/value.go�4type..hash.[2]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0780 type.int "".autotmp_0779 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[2]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�0type..eq.[2]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0784 ?"type.interface {} "".autotmp_0783 "type.interface {} "".autotmp_0782 _type.int "".autotmp_0781 Otype.int "".~r2  type.bool "".q *type.*[2]interface {} "".p  *type.*[2]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   @$GOROOT/src/go/constant/value.go�("".Value.ExactString �  �dH�%    H;avSH��H�Y H��tH�|$ H9;uH�#1�H�\$0H�\$8H�\$(H�$H�\$ H�[ ��H�L$H�D$H�L$0H�D$8H����    ��������
      �       �  0runtime.morestack_noctxt   @0  "".~r0  type.string ""..this  type."".Value 0N/ p 4p 
 G) Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�"".Value.Kind �  �dH�%    H;av=H��H�Y H��tH�|$H9;uH�#H�\$ H�$H�\$H�[(��H�\$H�\$(H����    ��������������
      v       �  0runtime.morestack_noctxt   0   "".~r0  type."".Kind ""..this  type."".Value  8 ` 6` 
 ;% Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�"".Value.String �  �dH�%    H;avSH��H�Y H��tH�|$ H9;uH�#1�H�\$0H�\$8H�\$(H�$H�\$ H�[0��H�L$H�D$H�L$0H�D$8H����    ��������
      �       �  0runtime.morestack_noctxt   @0  "".~r0  type.string ""..this  type."".Value 0N/ p 8p 
 G) Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�0"".Value.implementsValue �  �dH�%    H;av3H��H�Y H��tH�|$H9;uH�#H�\$H�$H�\$H�[8��H����    ��������
      v       �  0runtime.morestack_noctxt      ""..this  type."".Value . P :P 
 ; Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�0type..hash."".complexVal �  �dH�%    H;avmH��H�\$ H�$H�<$ tPH�\$(H�\$�    H�D$H�\$ H�$H�<$ t#H�$H�D$(H�D$�    H�\$H�\$0H��É%    �ԉ%    ��    �z�������������
      \  "runtime.interhash   �  "runtime.interhash   �  0runtime.morestack_noctxt   00  "".~r2  type.uintptr "".h type.uintptr "".p  &type.*"".complexVal 0V/0/ � � 
 -c Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�,type..eq."".complexVal �  �dH�%    H;a�  H��HH�\$XH�� ��   H�H�sH�\$PH�� ��   H�H�SH9���   H�D$(H�$H�T$0H�T$H�L$8H�L$H�t$@H�t$�    �\$ �� t}H�\$XH�� tnH�KH�sH�\$PH�� tWH�CH�SH9�u@H�D$(H�$H�T$0H�T$H�L$8H�L$H�t$@H�t$�    �\$ �� t
�D$`H��H��D$` H��HÉ륉��D$` H��HÉ�,���������    ��������������������
      �  runtime.ifaceeq   �  runtime.ifaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0791  type."".Value "".autotmp_0790  type."".Value "".autotmp_0789 ?type."".Value "".autotmp_0788 type."".Value "".~r2  type.bool "".q &type.*"".complexVal "".p  &type.*"".complexVal 8����	����� � �  s� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   @$GOROOT/src/go/constant/value.go�*"".(*complexVal).Kind �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�|$8 tH��   H�D$@H��0É%    ���    �V���������
      x  (go.string."constant"   �  ,go.string."complexVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  &type.*"".complexVal `_`	_ � <� 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�."".(*complexVal).String �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�t$8H�� t&H���    �    H�L$ H�D$(H�L$@H�D$HH��0É���    �7����������
      �  (go.string."constant"   �  ,go.string."complexVal"   �  $go.string."String"   �  "runtime.panicwrap   ��  runtime.duffcopy   �  ("".complexVal.String   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  &type.*"".complexVal `�_`_ � >�  �M Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�8"".(*complexVal).ExactString �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$@H�\$HH�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�t$8H�� t&H���    �    H�L$ H�D$(H�L$@H�D$HH��0É���    �7����������
      �  (go.string."constant"   �  ,go.string."complexVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   ��  runtime.duffcopy   �  2"".complexVal.ExactString   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  &type.*"".complexVal `�_`_ � @�  �M Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�@"".(*complexVal).implementsValue �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  ,go.string."complexVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  &type.*"".complexVal `s_`	_ � B� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�*"".(*unknownVal).Kind �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�|$8 t1�H�D$@H��0É%    ���    �[��������������
      x  (go.string."constant"   �  ,go.string."unknownVal"   �   go.string."Kind"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type."".Kind ""..this  &type.*"".unknownVal `z_`	_ � D� 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�."".(*unknownVal).String �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�|$8 t1�H�    H��   H�\$@H�D$HH��0É%    ���    �F���������
      |  (go.string."constant"   �  ,go.string."unknownVal"   �  $go.string."String"   �  "runtime.panicwrap   �  &go.string."unknown"   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  &type.*"".unknownVal `�_`	_ � F� 
 yG Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�8"".(*unknownVal).ExactString �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#1�H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�\$8H�� t!1�1�H�    H��   H�L$@H�D$HH��0É���    �F���������
      |  (go.string."constant"   �  ,go.string."unknownVal"   �  .go.string."ExactString"   �  "runtime.panicwrap   �  &go.string."unknown"   �  0runtime.morestack_noctxt   0`  "".~r0 type.string ""..this  &type.*"".unknownVal `�_`_ � H� 
 yG Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�@"".(*unknownVal).implementsValue �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$
   H�    H�\$ H�D$(   �    H�|$8 tH��0É%    ���    �b�����
      x  (go.string."constant"   �  ,go.string."unknownVal"   �  6go.string."implementsValue"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt   `  ""..this  &type.*"".unknownVal `s_`	_ � J� 
 w) Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�4type..hash.[3]interface {} �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  (runtime.nilinterhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_0796 type.int "".autotmp_0795 type.int "".~r2  type.uintptr "".h type.uintptr "".p  *type.*[3]interface {} PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   @$GOROOT/src/go/constant/value.go�0type..eq.[3]interface {} �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.efaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_0800 ?"type.interface {} "".autotmp_0799 "type.interface {} "".autotmp_0798 _type.int "".autotmp_0797 Otype.int "".~r2  type.bool "".q *type.*[3]interface {} "".p  *type.*[3]interface {} ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   @$GOROOT/src/go/constant/value.go�Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·d0110d631ecd4af0947009e36d46dc99             �.go.string.hdr."unknown"                       &go.string."unknown"   �&go.string."unknown"   unknown  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �(go.string.hdr."true"                        go.string."true"   � go.string."true"   
true  �*go.string.hdr."false"                       "go.string."false"   �"go.string."false"   false  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �&go.string.hdr."..."                       go.string."..."   �go.string."..."   ...  �Tgclocals·83ead081cd909acab0dcd88a450c1878                   �Tgclocals·f47057354ec566066f8688a4970cff5a                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �(go.string.hdr."%.6g"                        go.string."%.6g"   � go.string."%.6g"   
%.6g  �0go.string.hdr."%.6ge%+d"                       (go.string."%.6ge%+d"   �(go.string."%.6ge%+d"    %.6ge%+d  �Tgclocals·ec147618165580e6a5d760bf3329b6ac H  H             8           /   /   �Tgclocals·948c285cf1025b717e2658a3cccfd415 H  H                            �4go.string.hdr."(%s + %si)"             
          ,go.string."(%s + %si)"   �,go.string."(%s + %si)"    (%s + %si)  �Tgclocals·341b909b97472a89efab32cbd0761e34 (  (   	       �  �   �Tgclocals·23322ef3fd8702babe318da8c8d339e7 (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a19b4fb8a607611184c7491e4d9543cb 0  0          @   Py  Px   �Tgclocals·ae0b17ff166fa616635ce4bad0c70f06 0  0                   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·31b2ddfd7c7062d584469c95698a3e1d             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·5184031d3a32a42d85027f073f873668              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·b40f0f67eae216e69d0bb41a8427b144 (  (                 �Tgclocals·f7309186bf9eeb0f8ece2eb16f2dc110 (  (                �>8go.itab."".int64Val."".Value     �Tgclocals·4cf9735ef08c57d91ff7cf30faacc15b                   �Tgclocals·aa5118865dd28fc3eaacbfc830efb456                  �>4go.itab."".intVal."".Value     �Tgclocals·83ead081cd909acab0dcd88a450c1878                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �>4go.itab."".ratVal."".Value     �>8go.itab."".floatVal."".Value     �Tgclocals·549df0c0b9c1ff589e7323390661782b P  P                                �Tgclocals·add78ec634cef78099972ccd9d767bc6 P  P                               �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �><go.itab."".complexVal."".Value     �Tgclocals·4cf9735ef08c57d91ff7cf30faacc15b                   �Tgclocals·8c2f8f990ab0a90930a640c5478081b4                  �Tgclocals·e48b749e068cae7c3a399141c10fe5f0 (  (                 �Tgclocals·55cc6ee7528f0b48e5a6d9bfba36524a (  (                �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �><go.itab."".unknownVal."".Value     �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �>6go.itab."".boolVal."".Value     �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �>:go.itab."".stringVal."".Value     �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·f47057354ec566066f8688a4970cff5a                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·f56b2291fa344104975cb6587be42b9b                    �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·f56b2291fa344104975cb6587be42b9b                    ��go.string.hdr."MakeFromLiteral called with non-zero last argument"             2          |go.string."MakeFromLiteral called with non-zero last argument"   �|go.string."MakeFromLiteral called with non-zero last argument" p  fMakeFromLiteral called with non-zero last argument  �Ngo.string.hdr."%v is not a valid token"                       Fgo.string."%v is not a valid token"   �Fgo.string."%v is not a valid token" 0  0%v is not a valid token  �Tgclocals·e6d79eb2ebb897d590c99339e042c95b �  �	   ,                                          �                         �Tgclocals·03a89d916197104e2ad001cc20167921 X  X	                                  �:go.string.hdr."%v not a Bool"                       2go.string."%v not a Bool"   �2go.string."%v not a Bool"    %v not a Bool  �Tgclocals·60492e1505747e8ca36c9c8f244a1b59 8  8          �   0  0   0   �Tgclocals·aa52d274abdec77c8c6f0039727529fb 8  8                      �>go.string.hdr."%v not a String"                       6go.string."%v not a String"   �6go.string."%v not a String"     %v not a String  �Tgclocals·29c773ae5a332cdcf56287cee2ea280d 8  8            �  �   �   �Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc 8  8                      �:go.string.hdr."%v not an Int"                       2go.string."%v not an Int"   �2go.string."%v not an Int"    %v not an Int  �Tgclocals·1170e30e7a2c29fab9e9231402d8c543 @  @          �     a  a   a   �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·50c543803d8632f8d2f7062c2b1cdc18 @  @          �     a@  a   a   �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �<go.string.hdr."%v not a Float"                       4go.string."%v not a Float"   �4go.string."%v not a Float"    %v not a Float  �Tgclocals·82e7e0e6288447ba602a0db7dfa00c79 @  @               �!  �  �	   �Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 @  @                         �Tgclocals·82e7e0e6288447ba602a0db7dfa00c79 @  @               �!  �  �	   �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·9df74eb5f212c312a79ae7ef34903c32 @  @               �  �   �   �Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 @  @                         �<go.string.hdr."%v not numeric"                       4go.string."%v not numeric"   �4go.string."%v not numeric"    %v not numeric  �Tgclocals·8efb4299ccfc450a63c2e51c4c5be655 @  @             �! � �	  �Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 @  @                         �Tgclocals·305e11413380417cd9c7d2ae9b79dbaa H  H               �  �   �   �   �Tgclocals·47e744d05637aa546b45723fe9d2d977 H  H                            �Tgclocals·524aafe7d1228e5424d64f5d94771fbf                   �Tgclocals·3260b5c802f633fd6252c227878dd72a                  �Fgo.string.hdr."%v not Int or Float"                       >go.string."%v not Int or Float"   �>go.string."%v not Int or Float" 0  (%v not Int or Float  �Tgclocals·0000613cea0d43cb0624ba62b8fe2aca @  @               �  �   �   �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·c04ada1956856a77e3bc187a9e8a1dcc @  @               C       �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·5ff70dccce69b73e733742f8f6b97bd8 @  @                 C         �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·2bee6dd56e8b158e514a8950bd21767b 8  8          �� 0� 0� 0�  �Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc 8  8                      �Tgclocals·707962cf7cb527a8361df5d978b0d876 @  @           �  � �� �� ��  �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·5a22249a9b0f12f04d737839c0e5b8d8 @  @          � � � � �  �Tgclocals·a68b09a48716afad7ca7a02fe6add474 @  @                         �Tgclocals·9d7301afadfdafb7e149f098ce5d5791 8  8   
       �  �  �  �   �Tgclocals·ae09aea6c950f33bbc27842daf2e8ebc 8  8                      �Tgclocals·ba07643250a35734cb355a9fec6f55cc �  �   +           ` �     �     �     ��    �     �    �Tgclocals·1dbe3e1675327063a63a3ea108cf04bf H  H                            �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Xgo.string.hdr."invalid unary operation %s%v"                       Pgo.string."invalid unary operation %s%v"   �Pgo.string."invalid unary operation %s%v" @  :invalid unary operation %s%v  �Tgclocals·37508b3b9062b4dfe185a1b1456475c6 �  �   ,           x `�    x  �    y  �    x` �    x  �   | `�    |  �    ~  �    x  �/   x  �/   x ��/    �Tgclocals·33962f28c07936e169c43edefa5ca65b p  p                                           �6go.string.hdr."unreachable"                       .go.string."unreachable"   �.go.string."unreachable"    unreachable  �Tgclocals·e94709487fd39cb5e22f0477cb3700dd (  (                 �Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 (  (                �Tgclocals·6964cae77cc8ca448bf07954c3733ae6 �  �   P               �    ��   �   ��   � 0  ��   ��    ��   ��    ��   ��    ��   �    ���   �    ���  � 0  ���  ��    ��   �   ��   �   ��   �   ��   �/   ��   �   ��   �   ���  � �  ��   �/   ��   �   ��   �   ��   �   ��    �Tgclocals·7f2bc03eae9ababa8d2e476fa773c6e9 �  �                                                                         �bgo.string.hdr."invalid binary operation %v %s %v"             !          Zgo.string."invalid binary operation %v %s %v"   �Zgo.string."invalid binary operation %v %s %v" P  Dinvalid binary operation %v %s %v  �Tgclocals·bbced691e09928f29a52c25e48674f8c �  �'   \               8        � 8     `  � 8"      � 8"      � 8       � 9        � 9�       � :        � :�       � <        � <�       � 8 $      � 8$      � �        � 8@!      � 8!      � x        � 8       � 8      
 � 8        �? 8      � 8       � 8   � `� 8   � f� 8     f� 8    � � 8    �` � 8   � x� 8   �  x� 8   �g  � 8   f �� 8   `f �� 8    f �� 8 � ` �� 8 �     � 8       ���8        ��8     �  �� �Tgclocals·4dd66991891153e33d6808f41376a850 �  �'                                                                                                                            �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·8ead428b4183a0f1b19d8f59d3dde163             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·8ead428b4183a0f1b19d8f59d3dde163             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·8ead428b4183a0f1b19d8f59d3dde163             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·8ead428b4183a0f1b19d8f59d3dde163             �Lgo.string.hdr."invalid shift %v %s %d"                       Dgo.string."invalid shift %v %s %d"   �Dgo.string."invalid shift %v %s %d" 0  .invalid shift %v %s %d  �Tgclocals·4b6ac10bfefaa8263abce44bdd57d854 H  H          1         � � A�  �Tgclocals·0588ca1c52d0ec7f6ca12931a37dd289 H  H                            �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·f56b2291fa344104975cb6587be42b9b                    �Vgo.string.hdr."invalid comparison %v %s %v"                       Ngo.string."invalid comparison %v %s %v"   �Ngo.string."invalid comparison %v %s %v" @  8invalid comparison %v %s %v  �Tgclocals·5ea1f2fbb7a4500b5337d2bd0531ab03 �  �   '                1               '          �   �    ~    ~   A ~    �Tgclocals·8348f4c3fb43d484332abd834bc6b74d p  p                                           �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �<"".minInt64  $type.*math/big.Int   �<"".maxInt64  $type.*math/big.Int   �<"".floatVal0   type."".floatVal   �>"".initdone·  type.uint8   �*"".unknownVal.Kind·f              $"".unknownVal.Kind   �$"".boolVal.Kind·f              "".boolVal.Kind   �("".stringVal.Kind·f              """.stringVal.Kind   �&"".int64Val.Kind·f               "".int64Val.Kind   �""".intVal.Kind·f              "".intVal.Kind   �""".ratVal.Kind·f              "".ratVal.Kind   �&"".floatVal.Kind·f               "".floatVal.Kind   �*"".complexVal.Kind·f              $"".complexVal.Kind   �."".unknownVal.String·f              ("".unknownVal.String   �("".boolVal.String·f              """.boolVal.String   �,"".stringVal.String·f              &"".stringVal.String   �*"".int64Val.String·f              $"".int64Val.String   �&"".intVal.String·f               "".intVal.String   �&"".ratVal.String·f               "".ratVal.String   �*"".floatVal.String·f              $"".floatVal.String   �."".complexVal.String·f              ("".complexVal.String   �8"".unknownVal.ExactString·f              2"".unknownVal.ExactString   �2"".boolVal.ExactString·f              ,"".boolVal.ExactString   �6"".stringVal.ExactString·f              0"".stringVal.ExactString   �4"".int64Val.ExactString·f              ."".int64Val.ExactString   �0"".intVal.ExactString·f              *"".intVal.ExactString   �0"".ratVal.ExactString·f              *"".ratVal.ExactString   �4"".floatVal.ExactString·f              ."".floatVal.ExactString   �8"".complexVal.ExactString·f              2"".complexVal.ExactString   �@"".unknownVal.implementsValue·f              :"".unknownVal.implementsValue   �:"".boolVal.implementsValue·f              4"".boolVal.implementsValue   �>"".stringVal.implementsValue·f              8"".stringVal.implementsValue   �<"".int64Val.implementsValue·f              6"".int64Val.implementsValue   �8"".ratVal.implementsValue·f              2"".ratVal.implementsValue   �8"".intVal.implementsValue·f              2"".intVal.implementsValue   �<"".floatVal.implementsValue·f              6"".floatVal.implementsValue   �@"".complexVal.implementsValue·f              :"".complexVal.implementsValue   �"".newInt·f              "".newInt   �"".newRat·f              "".newRat   �"".newFloat·f              "".newFloat   �"".i64toi·f              "".i64toi   �"".i64tor·f              "".i64tor   �"".i64tof·f              "".i64tof   �"".itor·f              "".itor   �"".itof·f              "".itof   �"".rtof·f              "".rtof   �"".vtoc·f              "".vtoc   �"".makeInt·f              "".makeInt   �"".makeRat·f              "".makeRat   �"".makeFloat·f              "".makeFloat   �""".makeComplex·f              "".makeComplex   �4"".makeFloatFromLiteral·f              ."".makeFloatFromLiteral   �"".smallRat·f              "".smallRat   �""".MakeUnknown·f              "".MakeUnknown   �"".MakeBool·f              "".MakeBool   � "".MakeString·f              "".MakeString   �"".MakeInt64·f              "".MakeInt64   � "".MakeUint64·f              "".MakeUint64   �""".MakeFloat64·f              "".MakeFloat64   �*"".MakeFromLiteral·f              $"".MakeFromLiteral   �"".BoolVal·f              "".BoolVal   �"".StringVal·f              "".StringVal   �"".Int64Val·f              "".Int64Val   �"".Uint64Val·f              "".Uint64Val   � "".Float32Val·f              "".Float32Val   � "".Float64Val·f              "".Float64Val   �"".BitLen·f              "".BitLen   �"".Sign·f              "".Sign   �"".Bytes·f              "".Bytes   �&"".MakeFromBytes·f               "".MakeFromBytes   �"".Num·f              "".Num   �"".Denom·f              "".Denom   �"".MakeImag·f              "".MakeImag   �"".Real·f              "".Real   �"".Imag·f              "".Imag   �"".ToInt·f              "".ToInt   �"".ToFloat·f              "".ToFloat   �"".ToComplex·f              "".ToComplex   �"".is32bit·f              "".is32bit   �"".is63bit·f              "".is63bit   �"".UnaryOp·f              "".UnaryOp   �"".ord·f              "".ord   �"".match·f              "".match   �"".BinaryOp·f              "".BinaryOp   �"".add·f              "".add   �"".sub·f              "".sub   �"".mul·f              "".mul   �"".quo·f              "".quo   �"".Shift·f              "".Shift   �"".cmpZero·f              "".cmpZero   �"".Compare·f              "".Compare   �"".init·f              "".init   �"runtime.gcbits.01    �<go.string.hdr."*constant.Kind"                       4go.string."*constant.Kind"   �4go.string."*constant.Kind"    *constant.Kind  �type.*"".Kind  �  �              *��M 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."*constant.Kind"   p  ,go.weak.type.**"".Kind   �  type."".Kind   �runtime.gcbits.      �:go.string.hdr."constant.Kind"                       2go.string."constant.Kind"   �2go.string."constant.Kind"    constant.Kind  �(go.string.hdr."Kind"                        go.string."Kind"   � go.string."Kind"   
Kind  �6go.string.hdr."go/constant"                       .go.string."go/constant"   �.go.string."go/constant"    go/constant  �"go.importpath."".                       .go.string."go/constant"   �type."".Kind  �  �               �w�m �                                                                                0�  runtime.algarray   @  runtime.gcbits.   P  :go.string.hdr."constant.Kind"   p  type.*"".Kind   `� type."".Kind   �  (go.string.hdr."Kind"   �  "go.importpath."".   �� type."".Kind   �Bgo.string.hdr."*constant.boolVal"                       :go.string."*constant.boolVal"   �:go.string."*constant.boolVal" 0  $*constant.boolVal  �0go.string.hdr."constant"                       (go.string."constant"   �(go.string."constant"    constant  �.go.string.hdr."boolVal"                       &go.string."boolVal"   �&go.string."boolVal"   boolVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �,go.string.hdr."String"                       $go.string."String"   �$go.string."String"   String  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �6go.string.hdr."ExactString"                       .go.string."ExactString"   �.go.string."ExactString"    ExactString  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �>go.string.hdr."implementsValue"                       6go.string."implementsValue"   �6go.string."implementsValue"     implementsValue  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �\go.string.hdr."func(*constant.boolVal) string"                       Tgo.string."func(*constant.boolVal) string"   �Tgo.string."func(*constant.boolVal) string" @  >func(*constant.boolVal) string  �:type.func(*"".boolVal) string �  �              ��O 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(*constant.boolVal) string"   p  Lgo.weak.type.*func(*"".boolVal) string   �� :type.func(*"".boolVal) string   �� :type.func(*"".boolVal) string   �   type.*"".boolVal   �  type.string   ��go.typelink.func(*constant.boolVal) string	func(*"".boolVal) string              :type.func(*"".boolVal) string   �jgo.string.hdr."func(*constant.boolVal) constant.Kind"             %          bgo.string."func(*constant.boolVal) constant.Kind"   �bgo.string."func(*constant.boolVal) constant.Kind" P  Lfunc(*constant.boolVal) constant.Kind  �<type.func(*"".boolVal) "".Kind �  �              M�*� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(*constant.boolVal) constant.Kind"   p  Ngo.weak.type.*func(*"".boolVal) "".Kind   �� <type.func(*"".boolVal) "".Kind   �� <type.func(*"".boolVal) "".Kind   �   type.*"".boolVal   �  type."".Kind   ��go.typelink.func(*constant.boolVal) constant.Kind	func(*"".boolVal) "".Kind              <type.func(*"".boolVal) "".Kind   �Ngo.string.hdr."func(*constant.boolVal)"                       Fgo.string."func(*constant.boolVal)"   �Fgo.string."func(*constant.boolVal)" 0  0func(*constant.boolVal)  �,type.func(*"".boolVal) �  �              S� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."func(*constant.boolVal)"   p  >go.weak.type.*func(*"".boolVal)   �� ,type.func(*"".boolVal)   �� ,type.func(*"".boolVal)   �   type.*"".boolVal   �jgo.typelink.func(*constant.boolVal)	func(*"".boolVal)              ,type.func(*"".boolVal)   �:go.string.hdr."func() string"                       2go.string."func() string"   �2go.string."func() string"    func() string  �$type.func() string �  �              �m� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."func() string"   p  6go.weak.type.*func() string   �� $type.func() string   �� $type.func() string   �  type.string   �Ngo.typelink.func() string	func() string              $type.func() string   �Hgo.string.hdr."func() constant.Kind"                       @go.string."func() constant.Kind"   �@go.string."func() constant.Kind" 0  *func() constant.Kind  �&type.func() "".Kind �  �              N�h� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."func() constant.Kind"   p  8go.weak.type.*func() "".Kind   �� &type.func() "".Kind   �� &type.func() "".Kind   �  type."".Kind   �^go.typelink.func() constant.Kind	func() "".Kind              &type.func() "".Kind   �,go.string.hdr."func()"                       $go.string."func()"   �$go.string."func()"   func()  �type.func() �  �              ���� 3                                                                                                0�  runtime.algarray   @  "runtime.gcbits.01   P  ,go.string.hdr."func()"   p  (go.weak.type.*func()   �� type.func()   �� type.func()   �2go.typelink.func()	func()              type.func()   � type.*"".boolVal  �  �              �~3� 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."*constant.boolVal"   p  2go.weak.type.**"".boolVal   �  type."".boolVal   `�  type.*"".boolVal   ��  type.*"".boolVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  :type.func(*"".boolVal) string   �  2"".(*boolVal).ExactString   �  2"".(*boolVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  <type.func(*"".boolVal) "".Kind   �  $"".(*boolVal).Kind   �  $"".(*boolVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  :type.func(*"".boolVal) string   �  ("".(*boolVal).String   �  ("".(*boolVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  ,type.func(*"".boolVal)   �  :"".(*boolVal).implementsValue   �  :"".(*boolVal).implementsValue   �@go.string.hdr."constant.boolVal"                       8go.string."constant.boolVal"   �8go.string."constant.boolVal" 0  "constant.boolVal  �Zgo.string.hdr."func(constant.boolVal) string"                       Rgo.string."func(constant.boolVal) string"   �Rgo.string."func(constant.boolVal) string" @  <func(constant.boolVal) string  �8type.func("".boolVal) string �  �              )5� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."func(constant.boolVal) string"   p  Jgo.weak.type.*func("".boolVal) string   �� 8type.func("".boolVal) string   �� 8type.func("".boolVal) string   �  type."".boolVal   �  type.string   ��go.typelink.func(constant.boolVal) string	func("".boolVal) string              8type.func("".boolVal) string   �hgo.string.hdr."func(constant.boolVal) constant.Kind"             $          `go.string."func(constant.boolVal) constant.Kind"   �`go.string."func(constant.boolVal) constant.Kind" P  Jfunc(constant.boolVal) constant.Kind  �:type.func("".boolVal) "".Kind �  �               � 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  hgo.string.hdr."func(constant.boolVal) constant.Kind"   p  Lgo.weak.type.*func("".boolVal) "".Kind   �� :type.func("".boolVal) "".Kind   �� :type.func("".boolVal) "".Kind   �  type."".boolVal   �  type."".Kind   ��go.typelink.func(constant.boolVal) constant.Kind	func("".boolVal) "".Kind              :type.func("".boolVal) "".Kind   �Lgo.string.hdr."func(constant.boolVal)"                       Dgo.string."func(constant.boolVal)"   �Dgo.string."func(constant.boolVal)" 0  .func(constant.boolVal)  �*type.func("".boolVal) �  �              O; 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."func(constant.boolVal)"   p  <go.weak.type.*func("".boolVal)   �� *type.func("".boolVal)   �� *type.func("".boolVal)   �  type."".boolVal   �fgo.typelink.func(constant.boolVal)	func("".boolVal)              *type.func("".boolVal)   �type."".boolVal  �  �               ��
& �                                                                                                                                                                                                                                                                              :0@  runtime.algarray   @  runtime.gcbits.   P  @go.string.hdr."constant.boolVal"   p   type.*"".boolVal   `� type."".boolVal   �  .go.string.hdr."boolVal"   �  "go.importpath."".   �� type."".boolVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  8type.func("".boolVal) string   �  2"".(*boolVal).ExactString   �  ,"".boolVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  :type.func("".boolVal) "".Kind   �  $"".(*boolVal).Kind   �  "".boolVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  8type.func("".boolVal) string   �  ("".(*boolVal).String   �  """.boolVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  *type.func("".boolVal)   �  :"".(*boolVal).implementsValue   �  4"".boolVal.implementsValue   �Fgo.string.hdr."*constant.stringVal"                       >go.string."*constant.stringVal"   �>go.string."*constant.stringVal" 0  (*constant.stringVal  �2go.string.hdr."stringVal"             	          *go.string."stringVal"   �*go.string."stringVal"    stringVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �`go.string.hdr."func(*constant.stringVal) string"                        Xgo.string."func(*constant.stringVal) string"   �Xgo.string."func(*constant.stringVal) string" P  Bfunc(*constant.stringVal) string  �>type.func(*"".stringVal) string �  �              ��t� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(*constant.stringVal) string"   p  Pgo.weak.type.*func(*"".stringVal) string   �� >type.func(*"".stringVal) string   �� >type.func(*"".stringVal) string   �  $type.*"".stringVal   �  type.string   ��go.typelink.func(*constant.stringVal) string	func(*"".stringVal) string              >type.func(*"".stringVal) string   �ngo.string.hdr."func(*constant.stringVal) constant.Kind"             '          fgo.string."func(*constant.stringVal) constant.Kind"   �fgo.string."func(*constant.stringVal) constant.Kind" P  Pfunc(*constant.stringVal) constant.Kind  �@type.func(*"".stringVal) "".Kind �  �              �=�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ngo.string.hdr."func(*constant.stringVal) constant.Kind"   p  Rgo.weak.type.*func(*"".stringVal) "".Kind   �� @type.func(*"".stringVal) "".Kind   �� @type.func(*"".stringVal) "".Kind   �  $type.*"".stringVal   �  type."".Kind   ��go.typelink.func(*constant.stringVal) constant.Kind	func(*"".stringVal) "".Kind              @type.func(*"".stringVal) "".Kind   �Rgo.string.hdr."func(*constant.stringVal)"                       Jgo.string."func(*constant.stringVal)"   �Jgo.string."func(*constant.stringVal)" @  4func(*constant.stringVal)  �0type.func(*"".stringVal) �  �              ���� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func(*constant.stringVal)"   p  Bgo.weak.type.*func(*"".stringVal)   �� 0type.func(*"".stringVal)   �� 0type.func(*"".stringVal)   �  $type.*"".stringVal   �rgo.typelink.func(*constant.stringVal)	func(*"".stringVal)              0type.func(*"".stringVal)   �$type.*"".stringVal  �  �              ��Xf 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."*constant.stringVal"   p  6go.weak.type.**"".stringVal   �  "type."".stringVal   `� $type.*"".stringVal   �� $type.*"".stringVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  >type.func(*"".stringVal) string   �  6"".(*stringVal).ExactString   �  6"".(*stringVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  @type.func(*"".stringVal) "".Kind   �  ("".(*stringVal).Kind   �  ("".(*stringVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  >type.func(*"".stringVal) string   �  ,"".(*stringVal).String   �  ,"".(*stringVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  0type.func(*"".stringVal)   �  >"".(*stringVal).implementsValue   �  >"".(*stringVal).implementsValue   �Dgo.string.hdr."constant.stringVal"                       <go.string."constant.stringVal"   �<go.string."constant.stringVal" 0  &constant.stringVal  �^go.string.hdr."func(constant.stringVal) string"                       Vgo.string."func(constant.stringVal) string"   �Vgo.string."func(constant.stringVal) string" @  @func(constant.stringVal) string  �<type.func("".stringVal) string �  �              *F*� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(constant.stringVal) string"   p  Ngo.weak.type.*func("".stringVal) string   �� <type.func("".stringVal) string   �� <type.func("".stringVal) string   �  "type."".stringVal   �  type.string   ��go.typelink.func(constant.stringVal) string	func("".stringVal) string              <type.func("".stringVal) string   �lgo.string.hdr."func(constant.stringVal) constant.Kind"             &          dgo.string."func(constant.stringVal) constant.Kind"   �dgo.string."func(constant.stringVal) constant.Kind" P  Nfunc(constant.stringVal) constant.Kind  �>type.func("".stringVal) "".Kind �  �              ��		 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(constant.stringVal) constant.Kind"   p  Pgo.weak.type.*func("".stringVal) "".Kind   �� >type.func("".stringVal) "".Kind   �� >type.func("".stringVal) "".Kind   �  "type."".stringVal   �  type."".Kind   ��go.typelink.func(constant.stringVal) constant.Kind	func("".stringVal) "".Kind              >type.func("".stringVal) "".Kind   �Pgo.string.hdr."func(constant.stringVal)"                       Hgo.string."func(constant.stringVal)"   �Hgo.string."func(constant.stringVal)" @  2func(constant.stringVal)  �.type.func("".stringVal) �  �              :BC� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Pgo.string.hdr."func(constant.stringVal)"   p  @go.weak.type.*func("".stringVal)   �� .type.func("".stringVal)   �� .type.func("".stringVal)   �  "type."".stringVal   �ngo.typelink.func(constant.stringVal)	func("".stringVal)              .type.func("".stringVal)   �"type."".stringVal  �  �              �n�                                                                                                                                                                                                                                                                               :0�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."constant.stringVal"   p  $type.*"".stringVal   `� "type."".stringVal   �  2go.string.hdr."stringVal"   �  "go.importpath."".   �� "type."".stringVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  <type.func("".stringVal) string   �  6"".(*stringVal).ExactString   �  0"".stringVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  >type.func("".stringVal) "".Kind   �  ("".(*stringVal).Kind   �  """.stringVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  <type.func("".stringVal) string   �  ,"".(*stringVal).String   �  &"".stringVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  .type.func("".stringVal)   �  >"".(*stringVal).implementsValue   �  8"".stringVal.implementsValue   �Dgo.string.hdr."*constant.int64Val"                       <go.string."*constant.int64Val"   �<go.string."*constant.int64Val" 0  &*constant.int64Val  �0go.string.hdr."int64Val"                       (go.string."int64Val"   �(go.string."int64Val"    int64Val  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �^go.string.hdr."func(*constant.int64Val) string"                       Vgo.string."func(*constant.int64Val) string"   �Vgo.string."func(*constant.int64Val) string" @  @func(*constant.int64Val) string  �<type.func(*"".int64Val) string �  �              �֘ 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(*constant.int64Val) string"   p  Ngo.weak.type.*func(*"".int64Val) string   �� <type.func(*"".int64Val) string   �� <type.func(*"".int64Val) string   �  "type.*"".int64Val   �  type.string   ��go.typelink.func(*constant.int64Val) string	func(*"".int64Val) string              <type.func(*"".int64Val) string   �lgo.string.hdr."func(*constant.int64Val) constant.Kind"             &          dgo.string."func(*constant.int64Val) constant.Kind"   �dgo.string."func(*constant.int64Val) constant.Kind" P  Nfunc(*constant.int64Val) constant.Kind  �>type.func(*"".int64Val) "".Kind �  �              9 7 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(*constant.int64Val) constant.Kind"   p  Pgo.weak.type.*func(*"".int64Val) "".Kind   �� >type.func(*"".int64Val) "".Kind   �� >type.func(*"".int64Val) "".Kind   �  "type.*"".int64Val   �  type."".Kind   ��go.typelink.func(*constant.int64Val) constant.Kind	func(*"".int64Val) "".Kind              >type.func(*"".int64Val) "".Kind   �Pgo.string.hdr."func(*constant.int64Val)"                       Hgo.string."func(*constant.int64Val)"   �Hgo.string."func(*constant.int64Val)" @  2func(*constant.int64Val)  �.type.func(*"".int64Val) �  �              �k7w 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Pgo.string.hdr."func(*constant.int64Val)"   p  @go.weak.type.*func(*"".int64Val)   �� .type.func(*"".int64Val)   �� .type.func(*"".int64Val)   �  "type.*"".int64Val   �ngo.typelink.func(*constant.int64Val)	func(*"".int64Val)              .type.func(*"".int64Val)   �"type.*"".int64Val  �  �              ���� 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."*constant.int64Val"   p  4go.weak.type.**"".int64Val   �   type."".int64Val   `� "type.*"".int64Val   �� "type.*"".int64Val   �  6go.string.hdr."ExactString"   �  $type.func() string   �  <type.func(*"".int64Val) string   �  4"".(*int64Val).ExactString   �  4"".(*int64Val).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  >type.func(*"".int64Val) "".Kind   �  &"".(*int64Val).Kind   �  &"".(*int64Val).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  <type.func(*"".int64Val) string   �  *"".(*int64Val).String   �  *"".(*int64Val).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  .type.func(*"".int64Val)   �  <"".(*int64Val).implementsValue   �  <"".(*int64Val).implementsValue   �Bgo.string.hdr."constant.int64Val"                       :go.string."constant.int64Val"   �:go.string."constant.int64Val" 0  $constant.int64Val  �\go.string.hdr."func(constant.int64Val) string"                       Tgo.string."func(constant.int64Val) string"   �Tgo.string."func(constant.int64Val) string" @  >func(constant.int64Val) string  �:type.func("".int64Val) string �  �              �Yi� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(constant.int64Val) string"   p  Lgo.weak.type.*func("".int64Val) string   �� :type.func("".int64Val) string   �� :type.func("".int64Val) string   �   type."".int64Val   �  type.string   ��go.typelink.func(constant.int64Val) string	func("".int64Val) string              :type.func("".int64Val) string   �jgo.string.hdr."func(constant.int64Val) constant.Kind"             %          bgo.string."func(constant.int64Val) constant.Kind"   �bgo.string."func(constant.int64Val) constant.Kind" P  Lfunc(constant.int64Val) constant.Kind  �<type.func("".int64Val) "".Kind �  �              	}� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(constant.int64Val) constant.Kind"   p  Ngo.weak.type.*func("".int64Val) "".Kind   �� <type.func("".int64Val) "".Kind   �� <type.func("".int64Val) "".Kind   �   type."".int64Val   �  type."".Kind   ��go.typelink.func(constant.int64Val) constant.Kind	func("".int64Val) "".Kind              <type.func("".int64Val) "".Kind   �Ngo.string.hdr."func(constant.int64Val)"                       Fgo.string."func(constant.int64Val)"   �Fgo.string."func(constant.int64Val)" 0  0func(constant.int64Val)  �,type.func("".int64Val) �  �              ��Em 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."func(constant.int64Val)"   p  >go.weak.type.*func("".int64Val)   �� ,type.func("".int64Val)   �� ,type.func("".int64Val)   �   type."".int64Val   �jgo.typelink.func(constant.int64Val)	func("".int64Val)              ,type.func("".int64Val)   � type."".int64Val  �  �               �T �                                                                                                                                                                                                                                                                              :0�  runtime.algarray   @  runtime.gcbits.   P  Bgo.string.hdr."constant.int64Val"   p  "type.*"".int64Val   `�  type."".int64Val   �  0go.string.hdr."int64Val"   �  "go.importpath."".   ��  type."".int64Val   �  6go.string.hdr."ExactString"   �  $type.func() string   �  :type.func("".int64Val) string   �  4"".(*int64Val).ExactString   �  ."".int64Val.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  <type.func("".int64Val) "".Kind   �  &"".(*int64Val).Kind   �   "".int64Val.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  :type.func("".int64Val) string   �  *"".(*int64Val).String   �  $"".int64Val.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  ,type.func("".int64Val)   �  <"".(*int64Val).implementsValue   �  6"".int64Val.implementsValue   �@go.string.hdr."*constant.intVal"                       8go.string."*constant.intVal"   �8go.string."*constant.intVal" 0  "*constant.intVal  �,go.string.hdr."intVal"                       $go.string."intVal"   �$go.string."intVal"   intVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Zgo.string.hdr."func(*constant.intVal) string"                       Rgo.string."func(*constant.intVal) string"   �Rgo.string."func(*constant.intVal) string" @  <func(*constant.intVal) string  �8type.func(*"".intVal) string �  �              �L2 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."func(*constant.intVal) string"   p  Jgo.weak.type.*func(*"".intVal) string   �� 8type.func(*"".intVal) string   �� 8type.func(*"".intVal) string   �  type.*"".intVal   �  type.string   ��go.typelink.func(*constant.intVal) string	func(*"".intVal) string              8type.func(*"".intVal) string   �hgo.string.hdr."func(*constant.intVal) constant.Kind"             $          `go.string."func(*constant.intVal) constant.Kind"   �`go.string."func(*constant.intVal) constant.Kind" P  Jfunc(*constant.intVal) constant.Kind  �:type.func(*"".intVal) "".Kind �  �              �6C 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  hgo.string.hdr."func(*constant.intVal) constant.Kind"   p  Lgo.weak.type.*func(*"".intVal) "".Kind   �� :type.func(*"".intVal) "".Kind   �� :type.func(*"".intVal) "".Kind   �  type.*"".intVal   �  type."".Kind   ��go.typelink.func(*constant.intVal) constant.Kind	func(*"".intVal) "".Kind              :type.func(*"".intVal) "".Kind   �Lgo.string.hdr."func(*constant.intVal)"                       Dgo.string."func(*constant.intVal)"   �Dgo.string."func(*constant.intVal)" 0  .func(*constant.intVal)  �*type.func(*"".intVal) �  �              g+� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."func(*constant.intVal)"   p  <go.weak.type.*func(*"".intVal)   �� *type.func(*"".intVal)   �� *type.func(*"".intVal)   �  type.*"".intVal   �fgo.typelink.func(*constant.intVal)	func(*"".intVal)              *type.func(*"".intVal)   �type.*"".intVal  �  �              ���
 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*constant.intVal"   p  0go.weak.type.**"".intVal   �  type."".intVal   `� type.*"".intVal   �� type.*"".intVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  8type.func(*"".intVal) string   �  0"".(*intVal).ExactString   �  0"".(*intVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  :type.func(*"".intVal) "".Kind   �  """.(*intVal).Kind   �  """.(*intVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  8type.func(*"".intVal) string   �  &"".(*intVal).String   �  &"".(*intVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  *type.func(*"".intVal)   �  8"".(*intVal).implementsValue   �  8"".(*intVal).implementsValue   �>go.string.hdr."constant.intVal"                       6go.string."constant.intVal"   �6go.string."constant.intVal"     constant.intVal  �&go.string.hdr."val"                       go.string."val"   �go.string."val"   val  �Xgo.string.hdr."func(constant.intVal) string"                       Pgo.string."func(constant.intVal) string"   �Pgo.string."func(constant.intVal) string" @  :func(constant.intVal) string  �6type.func("".intVal) string �  �              �;�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."func(constant.intVal) string"   p  Hgo.weak.type.*func("".intVal) string   �� 6type.func("".intVal) string   �� 6type.func("".intVal) string   �  type."".intVal   �  type.string   �~go.typelink.func(constant.intVal) string	func("".intVal) string              6type.func("".intVal) string   �fgo.string.hdr."func(constant.intVal) constant.Kind"             #          ^go.string."func(constant.intVal) constant.Kind"   �^go.string."func(constant.intVal) constant.Kind" P  Hfunc(constant.intVal) constant.Kind  �8type.func("".intVal) "".Kind �  �              ��0 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(constant.intVal) constant.Kind"   p  Jgo.weak.type.*func("".intVal) "".Kind   �� 8type.func("".intVal) "".Kind   �� 8type.func("".intVal) "".Kind   �  type."".intVal   �  type."".Kind   ��go.typelink.func(constant.intVal) constant.Kind	func("".intVal) "".Kind              8type.func("".intVal) "".Kind   �Jgo.string.hdr."func(constant.intVal)"                       Bgo.string."func(constant.intVal)"   �Bgo.string."func(constant.intVal)" 0  ,func(constant.intVal)  �(type.func("".intVal) �  �               6D� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Jgo.string.hdr."func(constant.intVal)"   p  :go.weak.type.*func("".intVal)   �� (type.func("".intVal)   �� (type.func("".intVal)   �  type."".intVal   �bgo.typelink.func(constant.intVal)	func("".intVal)              (type.func("".intVal)   �type."".intVal  �  �              @��q 9                                                                                                                                                                                                                                                                                                                                            B0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."constant.intVal"   p  type.*"".intVal   �� type."".intVal   �  &go.string.hdr."val"   �  "go.importpath."".   �  $type.*math/big.Int   `� type."".intVal   �  ,go.string.hdr."intVal"   �  "go.importpath."".   �� type."".intVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  6type.func("".intVal) string   �  *"".intVal.ExactString   �  *"".intVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  8type.func("".intVal) "".Kind   �  "".intVal.Kind   �  "".intVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  6type.func("".intVal) string   �   "".intVal.String   �   "".intVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  (type.func("".intVal)   �  2"".intVal.implementsValue   �  2"".intVal.implementsValue   �@go.string.hdr."*constant.ratVal"                       8go.string."*constant.ratVal"   �8go.string."*constant.ratVal" 0  "*constant.ratVal  �,go.string.hdr."ratVal"                       $go.string."ratVal"   �$go.string."ratVal"   ratVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �Zgo.string.hdr."func(*constant.ratVal) string"                       Rgo.string."func(*constant.ratVal) string"   �Rgo.string."func(*constant.ratVal) string" @  <func(*constant.ratVal) string  �8type.func(*"".ratVal) string �  �              ��@ 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Zgo.string.hdr."func(*constant.ratVal) string"   p  Jgo.weak.type.*func(*"".ratVal) string   �� 8type.func(*"".ratVal) string   �� 8type.func(*"".ratVal) string   �  type.*"".ratVal   �  type.string   ��go.typelink.func(*constant.ratVal) string	func(*"".ratVal) string              8type.func(*"".ratVal) string   �hgo.string.hdr."func(*constant.ratVal) constant.Kind"             $          `go.string."func(*constant.ratVal) constant.Kind"   �`go.string."func(*constant.ratVal) constant.Kind" P  Jfunc(*constant.ratVal) constant.Kind  �:type.func(*"".ratVal) "".Kind �  �              ��/ 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  hgo.string.hdr."func(*constant.ratVal) constant.Kind"   p  Lgo.weak.type.*func(*"".ratVal) "".Kind   �� :type.func(*"".ratVal) "".Kind   �� :type.func(*"".ratVal) "".Kind   �  type.*"".ratVal   �  type."".Kind   ��go.typelink.func(*constant.ratVal) constant.Kind	func(*"".ratVal) "".Kind              :type.func(*"".ratVal) "".Kind   �Lgo.string.hdr."func(*constant.ratVal)"                       Dgo.string."func(*constant.ratVal)"   �Dgo.string."func(*constant.ratVal)" 0  .func(*constant.ratVal)  �*type.func(*"".ratVal) �  �              D�O 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."func(*constant.ratVal)"   p  <go.weak.type.*func(*"".ratVal)   �� *type.func(*"".ratVal)   �� *type.func(*"".ratVal)   �  type.*"".ratVal   �fgo.typelink.func(*constant.ratVal)	func(*"".ratVal)              *type.func(*"".ratVal)   �type.*"".ratVal  �  �              C'� 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*constant.ratVal"   p  0go.weak.type.**"".ratVal   �  type."".ratVal   `� type.*"".ratVal   �� type.*"".ratVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  8type.func(*"".ratVal) string   �  0"".(*ratVal).ExactString   �  0"".(*ratVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  :type.func(*"".ratVal) "".Kind   �  """.(*ratVal).Kind   �  """.(*ratVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  8type.func(*"".ratVal) string   �  &"".(*ratVal).String   �  &"".(*ratVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  *type.func(*"".ratVal)   �  8"".(*ratVal).implementsValue   �  8"".(*ratVal).implementsValue   �>go.string.hdr."constant.ratVal"                       6go.string."constant.ratVal"   �6go.string."constant.ratVal"     constant.ratVal  �Xgo.string.hdr."func(constant.ratVal) string"                       Pgo.string."func(constant.ratVal) string"   �Pgo.string."func(constant.ratVal) string" @  :func(constant.ratVal) string  �6type.func("".ratVal) string �  �              xti 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."func(constant.ratVal) string"   p  Hgo.weak.type.*func("".ratVal) string   �� 6type.func("".ratVal) string   �� 6type.func("".ratVal) string   �  type."".ratVal   �  type.string   �~go.typelink.func(constant.ratVal) string	func("".ratVal) string              6type.func("".ratVal) string   �fgo.string.hdr."func(constant.ratVal) constant.Kind"             #          ^go.string."func(constant.ratVal) constant.Kind"   �^go.string."func(constant.ratVal) constant.Kind" P  Hfunc(constant.ratVal) constant.Kind  �8type.func("".ratVal) "".Kind �  �              w��� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(constant.ratVal) constant.Kind"   p  Jgo.weak.type.*func("".ratVal) "".Kind   �� 8type.func("".ratVal) "".Kind   �� 8type.func("".ratVal) "".Kind   �  type."".ratVal   �  type."".Kind   ��go.typelink.func(constant.ratVal) constant.Kind	func("".ratVal) "".Kind              8type.func("".ratVal) "".Kind   �Jgo.string.hdr."func(constant.ratVal)"                       Bgo.string."func(constant.ratVal)"   �Bgo.string."func(constant.ratVal)" 0  ,func(constant.ratVal)  �(type.func("".ratVal) �  �              ��	� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Jgo.string.hdr."func(constant.ratVal)"   p  :go.weak.type.*func("".ratVal)   �� (type.func("".ratVal)   �� (type.func("".ratVal)   �  type."".ratVal   �bgo.typelink.func(constant.ratVal)	func("".ratVal)              (type.func("".ratVal)   �type."".ratVal  �  �              ��> 9                                                                                                                                                                                                                                                                                                                                            B0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."constant.ratVal"   p  type.*"".ratVal   �� type."".ratVal   �  &go.string.hdr."val"   �  "go.importpath."".   �  $type.*math/big.Rat   `� type."".ratVal   �  ,go.string.hdr."ratVal"   �  "go.importpath."".   �� type."".ratVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  6type.func("".ratVal) string   �  *"".ratVal.ExactString   �  *"".ratVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  8type.func("".ratVal) "".Kind   �  "".ratVal.Kind   �  "".ratVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  6type.func("".ratVal) string   �   "".ratVal.String   �   "".ratVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  (type.func("".ratVal)   �  2"".ratVal.implementsValue   �  2"".ratVal.implementsValue   �Dgo.string.hdr."*constant.floatVal"                       <go.string."*constant.floatVal"   �<go.string."*constant.floatVal" 0  &*constant.floatVal  �0go.string.hdr."floatVal"                       (go.string."floatVal"   �(go.string."floatVal"    floatVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �^go.string.hdr."func(*constant.floatVal) string"                       Vgo.string."func(*constant.floatVal) string"   �Vgo.string."func(*constant.floatVal) string" @  @func(*constant.floatVal) string  �<type.func(*"".floatVal) string �  �              \q]c 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(*constant.floatVal) string"   p  Ngo.weak.type.*func(*"".floatVal) string   �� <type.func(*"".floatVal) string   �� <type.func(*"".floatVal) string   �  "type.*"".floatVal   �  type.string   ��go.typelink.func(*constant.floatVal) string	func(*"".floatVal) string              <type.func(*"".floatVal) string   �lgo.string.hdr."func(*constant.floatVal) constant.Kind"             &          dgo.string."func(*constant.floatVal) constant.Kind"   �dgo.string."func(*constant.floatVal) constant.Kind" P  Nfunc(*constant.floatVal) constant.Kind  �>type.func(*"".floatVal) "".Kind �  �              xb�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(*constant.floatVal) constant.Kind"   p  Pgo.weak.type.*func(*"".floatVal) "".Kind   �� >type.func(*"".floatVal) "".Kind   �� >type.func(*"".floatVal) "".Kind   �  "type.*"".floatVal   �  type."".Kind   ��go.typelink.func(*constant.floatVal) constant.Kind	func(*"".floatVal) "".Kind              >type.func(*"".floatVal) "".Kind   �Pgo.string.hdr."func(*constant.floatVal)"                       Hgo.string."func(*constant.floatVal)"   �Hgo.string."func(*constant.floatVal)" @  2func(*constant.floatVal)  �.type.func(*"".floatVal) �  �              kґ 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Pgo.string.hdr."func(*constant.floatVal)"   p  @go.weak.type.*func(*"".floatVal)   �� .type.func(*"".floatVal)   �� .type.func(*"".floatVal)   �  "type.*"".floatVal   �ngo.typelink.func(*constant.floatVal)	func(*"".floatVal)              .type.func(*"".floatVal)   �"type.*"".floatVal  �  �              (�=k 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."*constant.floatVal"   p  4go.weak.type.**"".floatVal   �   type."".floatVal   `� "type.*"".floatVal   �� "type.*"".floatVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  <type.func(*"".floatVal) string   �  4"".(*floatVal).ExactString   �  4"".(*floatVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  >type.func(*"".floatVal) "".Kind   �  &"".(*floatVal).Kind   �  &"".(*floatVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  <type.func(*"".floatVal) string   �  *"".(*floatVal).String   �  *"".(*floatVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  .type.func(*"".floatVal)   �  <"".(*floatVal).implementsValue   �  <"".(*floatVal).implementsValue   �Bgo.string.hdr."constant.floatVal"                       :go.string."constant.floatVal"   �:go.string."constant.floatVal" 0  $constant.floatVal  �\go.string.hdr."func(constant.floatVal) string"                       Tgo.string."func(constant.floatVal) string"   �Tgo.string."func(constant.floatVal) string" @  >func(constant.floatVal) string  �:type.func("".floatVal) string �  �              ��P 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(constant.floatVal) string"   p  Lgo.weak.type.*func("".floatVal) string   �� :type.func("".floatVal) string   �� :type.func("".floatVal) string   �   type."".floatVal   �  type.string   ��go.typelink.func(constant.floatVal) string	func("".floatVal) string              :type.func("".floatVal) string   �jgo.string.hdr."func(constant.floatVal) constant.Kind"             %          bgo.string."func(constant.floatVal) constant.Kind"   �bgo.string."func(constant.floatVal) constant.Kind" P  Lfunc(constant.floatVal) constant.Kind  �<type.func("".floatVal) "".Kind �  �               wI| 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(constant.floatVal) constant.Kind"   p  Ngo.weak.type.*func("".floatVal) "".Kind   �� <type.func("".floatVal) "".Kind   �� <type.func("".floatVal) "".Kind   �   type."".floatVal   �  type."".Kind   ��go.typelink.func(constant.floatVal) constant.Kind	func("".floatVal) "".Kind              <type.func("".floatVal) "".Kind   �Ngo.string.hdr."func(constant.floatVal)"                       Fgo.string."func(constant.floatVal)"   �Fgo.string."func(constant.floatVal)" 0  0func(constant.floatVal)  �,type.func("".floatVal) �  �              �ֵ 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."func(constant.floatVal)"   p  >go.weak.type.*func("".floatVal)   �� ,type.func("".floatVal)   �� ,type.func("".floatVal)   �   type."".floatVal   �jgo.typelink.func(constant.floatVal)	func("".floatVal)              ,type.func("".floatVal)   � type."".floatVal  �  �              1�� 9                                                                                                                                                                                                                                                                                                                                            B0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."constant.floatVal"   p  "type.*"".floatVal   ��  type."".floatVal   �  &go.string.hdr."val"   �  "go.importpath."".   �  (type.*math/big.Float   `�  type."".floatVal   �  0go.string.hdr."floatVal"   �  "go.importpath."".   ��  type."".floatVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  :type.func("".floatVal) string   �  ."".floatVal.ExactString   �  ."".floatVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  <type.func("".floatVal) "".Kind   �   "".floatVal.Kind   �   "".floatVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  :type.func("".floatVal) string   �  $"".floatVal.String   �  $"".floatVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  ,type.func("".floatVal)   �  6"".floatVal.implementsValue   �  6"".floatVal.implementsValue   �"runtime.gcbits.03    �8go.string.hdr."interface {}"                       0go.string."interface {}"   �0go.string."interface {}"    interface {}  �"type.interface {} �  �              �W�                                                                 
0�  runtime.algarray   @  "runtime.gcbits.03   P  8go.string.hdr."interface {}"   p  4go.weak.type.*interface {}   �� "type.interface {}   �<go.string.hdr."[]interface {}"                       4go.string."[]interface {}"   �4go.string."[]interface {}"    []interface {}  �&type.[]interface {} �  �              p��/                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."[]interface {}"   p  8go.weak.type.*[]interface {}   �  "type.interface {}   �Rgo.typelink.[]interface {}	[]interface {}              &type.[]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[1]interface {}              4type..hash.[1]interface {}   �8type..eqfunc.[1]interface {}              0type..eq.[1]interface {}   �2type..alg.[1]interface {}                        <type..hashfunc.[1]interface {}     8type..eqfunc.[1]interface {}   �>go.string.hdr."[1]interface {}"                       6go.string."[1]interface {}"   �6go.string."[1]interface {}"     [1]interface {}  �(type.[1]interface {} �  �              P�[�                                                                0  2type..alg.[1]interface {}   @  "runtime.gcbits.03   P  >go.string.hdr."[1]interface {}"   p  :go.weak.type.*[1]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[1]interface {}	[1]interface {}              (type.[1]interface {}   �@go.string.hdr."*[1]interface {}"                       8go.string."*[1]interface {}"   �8go.string."*[1]interface {}" 0  "*[1]interface {}  �*type.*[1]interface {} �  �              ��5 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[1]interface {}"   p  <go.weak.type.**[1]interface {}   �  (type.[1]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[2]interface {}              4type..hash.[2]interface {}   �8type..eqfunc.[2]interface {}              0type..eq.[2]interface {}   �2type..alg.[2]interface {}                        <type..hashfunc.[2]interface {}     8type..eqfunc.[2]interface {}   �"runtime.gcbits.0f    �>go.string.hdr."[2]interface {}"                       6go.string."[2]interface {}"   �6go.string."[2]interface {}"     [2]interface {}  �(type.[2]interface {} �  �                ,Y��                                                                0  2type..alg.[2]interface {}   @  "runtime.gcbits.0f   P  >go.string.hdr."[2]interface {}"   p  :go.weak.type.*[2]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[2]interface {}	[2]interface {}              (type.[2]interface {}   �@go.string.hdr."*[2]interface {}"                       8go.string."*[2]interface {}"   �8go.string."*[2]interface {}" 0  "*[2]interface {}  �*type.*[2]interface {} �  �              �s-q 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[2]interface {}"   p  <go.weak.type.**[2]interface {}   �  (type.[2]interface {}   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6             �>go.string.hdr."*constant.Value"                       6go.string."*constant.Value"   �6go.string."*constant.Value"     *constant.Value  �type.*"".Value  �  �              ��7� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."*constant.Value"   p  .go.weak.type.**"".Value   �  type."".Value   �<go.string.hdr."constant.Value"                       4go.string."constant.Value"   �4go.string."constant.Value"    constant.Value  �*go.string.hdr."Value"                       "go.string."Value"   �"go.string."Value"   Value  �type."".Value  �  �              ׻9                                                                                                                                                                                                       $0�  runtime.algarray   @  "runtime.gcbits.03   P  <go.string.hdr."constant.Value"   p  type.*"".Value   �� type."".Value   �  6go.string.hdr."ExactString"   �  $type.func() string   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   `� type."".Value   �  *go.string.hdr."Value"   �  "go.importpath."".   �� type."".Value   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �8type..hashfunc."".complexVal              0type..hash."".complexVal   �4type..eqfunc."".complexVal              ,type..eq."".complexVal   �.type..alg."".complexVal                        8type..hashfunc."".complexVal     4type..eqfunc."".complexVal   �Hgo.string.hdr."*constant.complexVal"                       @go.string."*constant.complexVal"   �@go.string."*constant.complexVal" 0  **constant.complexVal  �4go.string.hdr."complexVal"             
          ,go.string."complexVal"   �,go.string."complexVal"    complexVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �bgo.string.hdr."func(*constant.complexVal) string"             !          Zgo.string."func(*constant.complexVal) string"   �Zgo.string."func(*constant.complexVal) string" P  Dfunc(*constant.complexVal) string  �@type.func(*"".complexVal) string �  �              <1W� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*constant.complexVal) string"   p  Rgo.weak.type.*func(*"".complexVal) string   �� @type.func(*"".complexVal) string   �� @type.func(*"".complexVal) string   �  &type.*"".complexVal   �  type.string   ��go.typelink.func(*constant.complexVal) string	func(*"".complexVal) string              @type.func(*"".complexVal) string   �pgo.string.hdr."func(*constant.complexVal) constant.Kind"             (          hgo.string."func(*constant.complexVal) constant.Kind"   �hgo.string."func(*constant.complexVal) constant.Kind" `  Rfunc(*constant.complexVal) constant.Kind  �Btype.func(*"".complexVal) "".Kind �  �              Ps= 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  pgo.string.hdr."func(*constant.complexVal) constant.Kind"   p  Tgo.weak.type.*func(*"".complexVal) "".Kind   �� Btype.func(*"".complexVal) "".Kind   �� Btype.func(*"".complexVal) "".Kind   �  &type.*"".complexVal   �  type."".Kind   ��go.typelink.func(*constant.complexVal) constant.Kind	func(*"".complexVal) "".Kind              Btype.func(*"".complexVal) "".Kind   �Tgo.string.hdr."func(*constant.complexVal)"                       Lgo.string."func(*constant.complexVal)"   �Lgo.string."func(*constant.complexVal)" @  6func(*constant.complexVal)  �2type.func(*"".complexVal) �  �              �4c 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Tgo.string.hdr."func(*constant.complexVal)"   p  Dgo.weak.type.*func(*"".complexVal)   �� 2type.func(*"".complexVal)   �� 2type.func(*"".complexVal)   �  &type.*"".complexVal   �vgo.typelink.func(*constant.complexVal)	func(*"".complexVal)              2type.func(*"".complexVal)   �&type.*"".complexVal  �  �              r�� 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."*constant.complexVal"   p  8go.weak.type.**"".complexVal   �  $type."".complexVal   `� &type.*"".complexVal   �� &type.*"".complexVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  @type.func(*"".complexVal) string   �  8"".(*complexVal).ExactString   �  8"".(*complexVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  Btype.func(*"".complexVal) "".Kind   �  *"".(*complexVal).Kind   �  *"".(*complexVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  @type.func(*"".complexVal) string   �  ."".(*complexVal).String   �  ."".(*complexVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  2type.func(*"".complexVal)   �  @"".(*complexVal).implementsValue   �  @"".(*complexVal).implementsValue   �Fgo.string.hdr."constant.complexVal"                       >go.string."constant.complexVal"   �>go.string."constant.complexVal" 0  (constant.complexVal  �$go.string.hdr."re"                       go.string."re"   �go.string."re"   re  �$go.string.hdr."im"                       go.string."im"   �go.string."im"   im  �`go.string.hdr."func(constant.complexVal) string"                        Xgo.string."func(constant.complexVal) string"   �Xgo.string."func(constant.complexVal) string" P  Bfunc(constant.complexVal) string  �>type.func("".complexVal) string �  �              gI	� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(constant.complexVal) string"   p  Pgo.weak.type.*func("".complexVal) string   �� >type.func("".complexVal) string   �� >type.func("".complexVal) string   �  $type."".complexVal   �  type.string   ��go.typelink.func(constant.complexVal) string	func("".complexVal) string              >type.func("".complexVal) string   �ngo.string.hdr."func(constant.complexVal) constant.Kind"             '          fgo.string."func(constant.complexVal) constant.Kind"   �fgo.string."func(constant.complexVal) constant.Kind" P  Pfunc(constant.complexVal) constant.Kind  �@type.func("".complexVal) "".Kind �  �              H�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ngo.string.hdr."func(constant.complexVal) constant.Kind"   p  Rgo.weak.type.*func("".complexVal) "".Kind   �� @type.func("".complexVal) "".Kind   �� @type.func("".complexVal) "".Kind   �  $type."".complexVal   �  type."".Kind   ��go.typelink.func(constant.complexVal) constant.Kind	func("".complexVal) "".Kind              @type.func("".complexVal) "".Kind   �Rgo.string.hdr."func(constant.complexVal)"                       Jgo.string."func(constant.complexVal)"   �Jgo.string."func(constant.complexVal)" @  4func(constant.complexVal)  �0type.func("".complexVal) �  �              ��� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func(constant.complexVal)"   p  Bgo.weak.type.*func("".complexVal)   �� 0type.func("".complexVal)   �� 0type.func("".complexVal)   �  $type."".complexVal   �rgo.typelink.func(constant.complexVal)	func("".complexVal)              0type.func("".complexVal)   �$type."".complexVal  �  �                �q��                                                                                                                                                                                                                                                                                                                                                                                    H0  .type..alg."".complexVal   @  "runtime.gcbits.0f   P  Fgo.string.hdr."constant.complexVal"   p  &type.*"".complexVal   �� $type."".complexVal   �  $go.string.hdr."re"   �  "go.importpath."".   �  type."".Value   �  $go.string.hdr."im"   �  "go.importpath."".   �  type."".Value   `� $type."".complexVal   �  4go.string.hdr."complexVal"   �  "go.importpath."".   �� $type."".complexVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  >type.func("".complexVal) string   �  8"".(*complexVal).ExactString   �  2"".complexVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  @type.func("".complexVal) "".Kind   �  *"".(*complexVal).Kind   �  $"".complexVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  >type.func("".complexVal) string   �  ."".(*complexVal).String   �  ("".complexVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  0type.func("".complexVal)   �  @"".(*complexVal).implementsValue   �  :"".complexVal.implementsValue   �Hgo.string.hdr."*constant.unknownVal"                       @go.string."*constant.unknownVal"   �@go.string."*constant.unknownVal" 0  **constant.unknownVal  �4go.string.hdr."unknownVal"             
          ,go.string."unknownVal"   �,go.string."unknownVal"    unknownVal  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·87d20ce1b58390b294df80b886db78bf             �bgo.string.hdr."func(*constant.unknownVal) string"             !          Zgo.string."func(*constant.unknownVal) string"   �Zgo.string."func(*constant.unknownVal) string" P  Dfunc(*constant.unknownVal) string  �@type.func(*"".unknownVal) string �  �              �� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*constant.unknownVal) string"   p  Rgo.weak.type.*func(*"".unknownVal) string   �� @type.func(*"".unknownVal) string   �� @type.func(*"".unknownVal) string   �  &type.*"".unknownVal   �  type.string   ��go.typelink.func(*constant.unknownVal) string	func(*"".unknownVal) string              @type.func(*"".unknownVal) string   �pgo.string.hdr."func(*constant.unknownVal) constant.Kind"             (          hgo.string."func(*constant.unknownVal) constant.Kind"   �hgo.string."func(*constant.unknownVal) constant.Kind" `  Rfunc(*constant.unknownVal) constant.Kind  �Btype.func(*"".unknownVal) "".Kind �  �              3��@ 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  pgo.string.hdr."func(*constant.unknownVal) constant.Kind"   p  Tgo.weak.type.*func(*"".unknownVal) "".Kind   �� Btype.func(*"".unknownVal) "".Kind   �� Btype.func(*"".unknownVal) "".Kind   �  &type.*"".unknownVal   �  type."".Kind   ��go.typelink.func(*constant.unknownVal) constant.Kind	func(*"".unknownVal) "".Kind              Btype.func(*"".unknownVal) "".Kind   �Tgo.string.hdr."func(*constant.unknownVal)"                       Lgo.string."func(*constant.unknownVal)"   �Lgo.string."func(*constant.unknownVal)" @  6func(*constant.unknownVal)  �2type.func(*"".unknownVal) �  �              ?k� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Tgo.string.hdr."func(*constant.unknownVal)"   p  Dgo.weak.type.*func(*"".unknownVal)   �� 2type.func(*"".unknownVal)   �� 2type.func(*"".unknownVal)   �  &type.*"".unknownVal   �vgo.typelink.func(*constant.unknownVal)	func(*"".unknownVal)              2type.func(*"".unknownVal)   �&type.*"".unknownVal  �  �              �݈) 6                                                                                                                                                                                                                                                                                      80�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."*constant.unknownVal"   p  8go.weak.type.**"".unknownVal   �  $type."".unknownVal   `� &type.*"".unknownVal   �� &type.*"".unknownVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  @type.func(*"".unknownVal) string   �  8"".(*unknownVal).ExactString   �  8"".(*unknownVal).ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  Btype.func(*"".unknownVal) "".Kind   �  *"".(*unknownVal).Kind   �  *"".(*unknownVal).Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  @type.func(*"".unknownVal) string   �  ."".(*unknownVal).String   �  ."".(*unknownVal).String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  2type.func(*"".unknownVal)   �  @"".(*unknownVal).implementsValue   �  @"".(*unknownVal).implementsValue   �Fgo.string.hdr."constant.unknownVal"                       >go.string."constant.unknownVal"   �>go.string."constant.unknownVal" 0  (constant.unknownVal  �`go.string.hdr."func(constant.unknownVal) string"                        Xgo.string."func(constant.unknownVal) string"   �Xgo.string."func(constant.unknownVal) string" P  Bfunc(constant.unknownVal) string  �>type.func("".unknownVal) string �  �              :�hL 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(constant.unknownVal) string"   p  Pgo.weak.type.*func("".unknownVal) string   �� >type.func("".unknownVal) string   �� >type.func("".unknownVal) string   �  $type."".unknownVal   �  type.string   ��go.typelink.func(constant.unknownVal) string	func("".unknownVal) string              >type.func("".unknownVal) string   �ngo.string.hdr."func(constant.unknownVal) constant.Kind"             '          fgo.string."func(constant.unknownVal) constant.Kind"   �fgo.string."func(constant.unknownVal) constant.Kind" P  Pfunc(constant.unknownVal) constant.Kind  �@type.func("".unknownVal) "".Kind �  �              ��
{ 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ngo.string.hdr."func(constant.unknownVal) constant.Kind"   p  Rgo.weak.type.*func("".unknownVal) "".Kind   �� @type.func("".unknownVal) "".Kind   �� @type.func("".unknownVal) "".Kind   �  $type."".unknownVal   �  type."".Kind   ��go.typelink.func(constant.unknownVal) constant.Kind	func("".unknownVal) "".Kind              @type.func("".unknownVal) "".Kind   �Rgo.string.hdr."func(constant.unknownVal)"                       Jgo.string."func(constant.unknownVal)"   �Jgo.string."func(constant.unknownVal)" @  4func(constant.unknownVal)  �0type.func("".unknownVal) �  �              ���v 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func(constant.unknownVal)"   p  Bgo.weak.type.*func("".unknownVal)   �� 0type.func("".unknownVal)   �� 0type.func("".unknownVal)   �  $type."".unknownVal   �rgo.typelink.func(constant.unknownVal)	func("".unknownVal)              0type.func("".unknownVal)   �$type."".unknownVal  �  �                �|~? �                                                                                                                                                                                                                                                                                                      <0   runtime.algarray   @  runtime.gcbits.   P  Fgo.string.hdr."constant.unknownVal"   p  &type.*"".unknownVal   �� $type."".unknownVal   `� $type."".unknownVal   �  4go.string.hdr."unknownVal"   �  "go.importpath."".   �� $type."".unknownVal   �  6go.string.hdr."ExactString"   �  $type.func() string   �  >type.func("".unknownVal) string   �  8"".(*unknownVal).ExactString   �  2"".unknownVal.ExactString   �  (go.string.hdr."Kind"   �  &type.func() "".Kind   �  @type.func("".unknownVal) "".Kind   �  *"".(*unknownVal).Kind   �  $"".unknownVal.Kind   �  ,go.string.hdr."String"   �  $type.func() string   �  >type.func("".unknownVal) string   �  ."".(*unknownVal).String   �  ("".unknownVal.String   �  >go.string.hdr."implementsValue"   �  "go.importpath."".   �  type.func()   �  0type.func("".unknownVal)   �  @"".(*unknownVal).implementsValue   �  :"".unknownVal.implementsValue   �.go.string.hdr."[]uint8"                       &go.string."[]uint8"   �&go.string."[]uint8"   []uint8  �type.[]uint8 �  �              �~.8                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  .go.string.hdr."[]uint8"   p  *go.weak.type.*[]uint8   �  type.uint8   �6go.typelink.[]uint8	[]uint8              type.[]uint8   �4go.string.hdr."[]big.Word"             
          ,go.string."[]big.Word"   �,go.string."[]big.Word"    []big.Word  �(type.[]math/big.Word �  �              =ҌN                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."[]big.Word"   p  :go.weak.type.*[]math/big.Word   �  $type.math/big.Word   �Lgo.typelink.[]big.Word	[]math/big.Word              (type.[]math/big.Word   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �<type..hashfunc.[3]interface {}              4type..hash.[3]interface {}   �8type..eqfunc.[3]interface {}              0type..eq.[3]interface {}   �2type..alg.[3]interface {}                        <type..hashfunc.[3]interface {}     8type..eqfunc.[3]interface {}   �"runtime.gcbits.3f   ? �>go.string.hdr."[3]interface {}"                       6go.string."[3]interface {}"   �6go.string."[3]interface {}"     [3]interface {}  �(type.[3]interface {} �  �0       0       ���                                                                0  2type..alg.[3]interface {}   @  "runtime.gcbits.3f   P  >go.string.hdr."[3]interface {}"   p  :go.weak.type.*[3]interface {}   �  "type.interface {}   �  &type.[]interface {}   �Vgo.typelink.[3]interface {}	[3]interface {}              (type.[3]interface {}   �@go.string.hdr."*[3]interface {}"                       8go.string."*[3]interface {}"   �8go.string."*[3]interface {}" 0  "*[3]interface {}  �*type.*[3]interface {} �  �              ��� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*[3]interface {}"   p  <go.weak.type.**[3]interface {}   �  (type.[3]interface {}   �&go.string.hdr."fmt"                       go.string."fmt"   �go.string."fmt"   fmt  �$go.importpath.fmt.                       go.string."fmt"   �(go.string.hdr."math"                        go.string."math"   � go.string."math"   
math  �&go.importpath.math.                        go.string."math"   �.go.string.hdr."strconv"                       &go.string."strconv"   �&go.string."strconv"   strconv  �,go.importpath.strconv.                       &go.string."strconv"   �8go.string.hdr."unicode/utf8"                       0go.string."unicode/utf8"   �0go.string."unicode/utf8"    unicode/utf8  �6go.importpath.unicode/utf8.                       0go.string."unicode/utf8"   �0go.string.hdr."go/token"                       (go.string."go/token"   �(go.string."go/token"    go/token  �.go.importpath.go/token.                       (go.string."go/token"   �0go.string.hdr."math/big"                       (go.string."math/big"   �(go.string."math/big"    math/big  �.go.importpath.math/big.                       (go.string."math/big"   �*"".(*boolVal).Kind·f              $"".(*boolVal).Kind   �."".(*boolVal).String·f              ("".(*boolVal).String   �8"".(*boolVal).ExactString·f              2"".(*boolVal).ExactString   �@"".(*boolVal).implementsValue·f              :"".(*boolVal).implementsValue   �."".(*stringVal).Kind·f              ("".(*stringVal).Kind   �2"".(*stringVal).String·f              ,"".(*stringVal).String   �<"".(*stringVal).ExactString·f              6"".(*stringVal).ExactString   �D"".(*stringVal).implementsValue·f              >"".(*stringVal).implementsValue   �,"".(*int64Val).Kind·f              &"".(*int64Val).Kind   �0"".(*int64Val).String·f              *"".(*int64Val).String   �:"".(*int64Val).ExactString·f              4"".(*int64Val).ExactString   �B"".(*int64Val).implementsValue·f              <"".(*int64Val).implementsValue   �("".(*intVal).Kind·f              """.(*intVal).Kind   �,"".(*intVal).String·f              &"".(*intVal).String   �6"".(*intVal).ExactString·f              0"".(*intVal).ExactString   �>"".(*intVal).implementsValue·f              8"".(*intVal).implementsValue   �("".(*ratVal).Kind·f              """.(*ratVal).Kind   �,"".(*ratVal).String·f              &"".(*ratVal).String   �6"".(*ratVal).ExactString·f              0"".(*ratVal).ExactString   �>"".(*ratVal).implementsValue·f              8"".(*ratVal).implementsValue   �,"".(*floatVal).Kind·f              &"".(*floatVal).Kind   �0"".(*floatVal).String·f              *"".(*floatVal).String   �:"".(*floatVal).ExactString·f              4"".(*floatVal).ExactString   �B"".(*floatVal).implementsValue·f              <"".(*floatVal).implementsValue   �:type..hash.[1]interface {}·f              4type..hash.[1]interface {}   �6type..eq.[1]interface {}·f              0type..eq.[1]interface {}   �:type..hash.[2]interface {}·f              4type..hash.[2]interface {}   �6type..eq.[2]interface {}·f              0type..eq.[2]interface {}   �."".Value.ExactString·f              ("".Value.ExactString   � "".Value.Kind·f              "".Value.Kind   �$"".Value.String·f              "".Value.String   �6"".Value.implementsValue·f              0"".Value.implementsValue   �6type..hash."".complexVal·f              0type..hash."".complexVal   �2type..eq."".complexVal·f              ,type..eq."".complexVal   �0"".(*complexVal).Kind·f              *"".(*complexVal).Kind   �4"".(*complexVal).String·f              ."".(*complexVal).String   �>"".(*complexVal).ExactString·f              8"".(*complexVal).ExactString   �F"".(*complexVal).implementsValue·f              @"".(*complexVal).implementsValue   �0"".(*unknownVal).Kind·f              *"".(*unknownVal).Kind   �4"".(*unknownVal).String·f              ."".(*unknownVal).String   �>"".(*unknownVal).ExactString·f              8"".(*unknownVal).ExactString   �F"".(*unknownVal).implementsValue·f              @"".(*unknownVal).implementsValue   �:type..hash.[3]interface {}·f              4type..hash.[3]interface {}   �6type..eq.[3]interface {}·f              0type..eq.[3]interface {}   ��go13ld                                                                                                                                                                                  usr/local/go/pkg/linux_amd64/go/doc.a                                                               0100644 0000000 0000000 00001554554 13101127332 016020  0                                                                                                    ustar 00                                                                0000000 0000000                                                                                                                                                                        !<arch>
__.PKGDEF       0           0     0     644     9966      `
go object linux amd64 go1.6.4 X:none
build id "08f71260798a3e1fddbdd2322479689e06f7f5a2"

$$
package doc
	import io "io"
	import regexp "regexp"
	import unicode "unicode"
	import sort "sort"
	import strings "strings"
	import utf8 "unicode/utf8"
	import strconv "strconv"
	import template "text/template"
	import ast "go/ast"
	import token "go/token"
	import path "path"
	type @"io".Writer interface { Write(@"io".p []byte) (@"io".n int, @"io".err error) }
	func @"".ToHTML (@"".w·1 @"io".Writer, @"".text·2 string, @"".words·3 map[string]string "esc:0x1")
	func @"".ToText (@"".w·1 @"io".Writer, @"".text·2 string, @"".indent·3 string, @"".preIndent·4 string "esc:0x1", @"".width·5 int)
	type @"go/token".Pos int
	func (@"go/token".p·2 @"go/token".Pos) IsValid () (? bool) { return @"go/token".p·2 != @"go/token".Pos(0x0) }
	type @"".Note struct { Pos @"go/token".Pos; End @"go/token".Pos; UID string; Body string }
	type @"go/ast".Comment struct { Slash @"go/token".Pos; Text string }
	func (@"go/ast".c·2 *@"go/ast".Comment "esc:0x1") End () (? @"go/token".Pos) { return @"go/token".Pos(int(@"go/ast".c·2.Slash) + len(@"go/ast".c·2.Text)) }
	func (@"go/ast".c·2 *@"go/ast".Comment "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".c·2.Slash }
	type @"go/ast".CommentGroup struct { List []*@"go/ast".Comment }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x1") End () (? @"go/token".Pos) { return @"go/ast".g·2.List[len(@"go/ast".g·2.List) - int(0x1)].End() }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".g·2.List[int(0x0)].Pos() }
	func (@"go/ast".g·2 *@"go/ast".CommentGroup "esc:0x9") Text () (? string)
	type @"go/token".Token int
	func (@"go/token".tok·2 @"go/token".Token) IsKeyword () (? bool) { return @"go/token".Token(0x3c) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0x56) }
	func (@"go/token".tok·2 @"go/token".Token) IsLiteral () (? bool) { return @"go/token".Token(0x3) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0xa) }
	func (@"go/token".tok·2 @"go/token".Token) IsOperator () (? bool) { return @"go/token".Token(0xb) < @"go/token".tok·2 && @"go/token".tok·2 < @"go/token".Token(0x3b) }
	func (@"go/token".op·2 @"go/token".Token) Precedence () (? int)
	func (@"go/token".tok·2 @"go/token".Token) String () (? string)
	type @"go/ast".Spec interface { End() (? @"go/token".Pos); Pos() (? @"go/token".Pos); @"go/ast".specNode() }
	type @"go/ast".GenDecl struct { Doc *@"go/ast".CommentGroup; TokPos @"go/token".Pos; Tok @"go/token".Token; Lparen @"go/token".Pos; Specs []@"go/ast".Spec; Rparen @"go/token".Pos }
	func (@"go/ast".d·2 *@"go/ast".GenDecl "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".d·2 *@"go/ast".GenDecl "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".d·2.TokPos }
	func (? *@"go/ast".GenDecl) @"go/ast".declNode () {  }
	type @"".Value struct { Doc string; Names []string; Decl *@"go/ast".GenDecl; @"".order int }
	type @"go/ast".ObjKind int
	func (@"go/ast".kind·2 @"go/ast".ObjKind) String () (? string) { return @"go/ast".objKindStrings[@"go/ast".kind·2] }
	type @"go/ast".Object struct { Kind @"go/ast".ObjKind; Name string; Decl interface {}; Data interface {}; Type interface {} }
	func (@"go/ast".obj·2 *@"go/ast".Object "esc:0x1") Pos () (? @"go/token".Pos)
	type @"go/ast".Ident struct { NamePos @"go/token".Pos; Name string; Obj *@"go/ast".Object }
	func (@"go/ast".x·2 *@"go/ast".Ident "esc:0x1") End () (? @"go/token".Pos) { return @"go/token".Pos(int(@"go/ast".x·2.NamePos) + len(@"go/ast".x·2.Name)) }
	func (@"go/ast".id·2 *@"go/ast".Ident "esc:0x1") IsExported () (? bool)
	func (@"go/ast".x·2 *@"go/ast".Ident "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".x·2.NamePos }
	func (@"go/ast".id·2 *@"go/ast".Ident "esc:0x22") String () (? string) { if @"go/ast".id·2 != nil { return @"go/ast".id·2.Name }; return string("<nil>") }
	func (? *@"go/ast".Ident) @"go/ast".exprNode () {  }
	type @"go/ast".Expr interface { End() (? @"go/token".Pos); Pos() (? @"go/token".Pos); @"go/ast".exprNode() }
	type @"go/ast".BasicLit struct { ValuePos @"go/token".Pos; Kind @"go/token".Token; Value string }
	func (@"go/ast".x·2 *@"go/ast".BasicLit "esc:0x1") End () (? @"go/token".Pos) { return @"go/token".Pos(int(@"go/ast".x·2.ValuePos) + len(@"go/ast".x·2.Value)) }
	func (@"go/ast".x·2 *@"go/ast".BasicLit "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".x·2.ValuePos }
	func (? *@"go/ast".BasicLit) @"go/ast".exprNode () {  }
	type @"go/ast".Field struct { Doc *@"go/ast".CommentGroup; Names []*@"go/ast".Ident; Type @"go/ast".Expr; Tag *@"go/ast".BasicLit; Comment *@"go/ast".CommentGroup }
	func (@"go/ast".f·2 *@"go/ast".Field "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".f·2 *@"go/ast".Field "esc:0x9") Pos () (? @"go/token".Pos)
	type @"go/ast".FieldList struct { Opening @"go/token".Pos; List []*@"go/ast".Field; Closing @"go/token".Pos }
	func (@"go/ast".f·2 *@"go/ast".FieldList "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".f·2 *@"go/ast".FieldList "esc:0x1") NumFields () (? int)
	func (@"go/ast".f·2 *@"go/ast".FieldList "esc:0x9") Pos () (? @"go/token".Pos)
	type @"go/ast".FuncType struct { Func @"go/token".Pos; Params *@"go/ast".FieldList; Results *@"go/ast".FieldList }
	func (@"go/ast".x·2 *@"go/ast".FuncType "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".x·2 *@"go/ast".FuncType "esc:0x9") Pos () (? @"go/token".Pos)
	func (? *@"go/ast".FuncType) @"go/ast".exprNode () {  }
	type @"go/ast".Stmt interface { End() (? @"go/token".Pos); Pos() (? @"go/token".Pos); @"go/ast".stmtNode() }
	type @"go/ast".BlockStmt struct { Lbrace @"go/token".Pos; List []@"go/ast".Stmt; Rbrace @"go/token".Pos }
	func (@"go/ast".s·2 *@"go/ast".BlockStmt "esc:0x1") End () (? @"go/token".Pos) { return @"go/ast".s·2.Rbrace + @"go/token".Pos(0x1) }
	func (@"go/ast".s·2 *@"go/ast".BlockStmt "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".s·2.Lbrace }
	func (? *@"go/ast".BlockStmt) @"go/ast".stmtNode () {  }
	type @"go/ast".FuncDecl struct { Doc *@"go/ast".CommentGroup; Recv *@"go/ast".FieldList; Name *@"go/ast".Ident; Type *@"go/ast".FuncType; Body *@"go/ast".BlockStmt }
	func (@"go/ast".d·2 *@"go/ast".FuncDecl "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".d·2 *@"go/ast".FuncDecl "esc:0x9") Pos () (? @"go/token".Pos)
	func (? *@"go/ast".FuncDecl) @"go/ast".declNode () {  }
	type @"".Func struct { Doc string; Name string; Decl *@"go/ast".FuncDecl; Recv string; Orig string; Level int }
	type @"".Type struct { Doc string; Name string; Decl *@"go/ast".GenDecl; Consts []*@"".Value; Vars []*@"".Value; Funcs []*@"".Func; Methods []*@"".Func }
	type @"".Filter func(? string) (? bool)
	type @"".Package struct { Doc string; Name string; ImportPath string; Imports []string; Filenames []string; Notes map[string][]*@"".Note; Bugs []string; Consts []*@"".Value; Types []*@"".Type; Vars []*@"".Value; Funcs []*@"".Func }
	func (@"".p·1 *@"".Package "esc:0x9") Filter (@"".f·2 @"".Filter "esc:0x1")
	type @"".Mode int
	const @"".AllDecls @"".Mode = 0x1
	const @"".AllMethods @"".Mode = 0x2
	type @"go/ast".Scope struct { Outer *@"go/ast".Scope; Objects map[string]*@"go/ast".Object }
	func (@"go/ast".s·2 *@"go/ast".Scope "esc:0x1") Insert (@"go/ast".obj·3 *@"go/ast".Object) (@"go/ast".alt·1 *@"go/ast".Object) { if @"go/ast".alt·1 = @"go/ast".s·2.Objects[@"go/ast".obj·3.Name]; @"go/ast".alt·1 == nil { @"go/ast".s·2.Objects[@"go/ast".obj·3.Name] = @"go/ast".obj·3 }; return  }
	func (@"go/ast".s·2 *@"go/ast".Scope "esc:0x1") Lookup (@"go/ast".name·3 string "esc:0x1") (? *@"go/ast".Object) { return @"go/ast".s·2.Objects[@"go/ast".name·3] }
	func (@"go/ast".s·2 *@"go/ast".Scope) String () (? string)
	type @"go/ast".Decl interface { End() (? @"go/token".Pos); Pos() (? @"go/token".Pos); @"go/ast".declNode() }
	type @"go/ast".ImportSpec struct { Doc *@"go/ast".CommentGroup; Name *@"go/ast".Ident; Path *@"go/ast".BasicLit; Comment *@"go/ast".CommentGroup; EndPos @"go/token".Pos }
	func (@"go/ast".s·2 *@"go/ast".ImportSpec "esc:0x1") End () (? @"go/token".Pos) { if @"go/ast".s·2.EndPos != @"go/token".Pos(0x0) { return @"go/ast".s·2.EndPos }; return @"go/ast".s·2.Path.End() }
	func (@"go/ast".s·2 *@"go/ast".ImportSpec "esc:0x1") Pos () (? @"go/token".Pos) { if @"go/ast".s·2.Name != nil { return @"go/ast".s·2.Name.Pos() }; return @"go/ast".s·2.Path.Pos() }
	func (? *@"go/ast".ImportSpec) @"go/ast".specNode () {  }
	type @"go/ast".File struct { Doc *@"go/ast".CommentGroup; Package @"go/token".Pos; Name *@"go/ast".Ident; Decls []@"go/ast".Decl; Scope *@"go/ast".Scope; Imports []*@"go/ast".ImportSpec; Unresolved []*@"go/ast".Ident; Comments []*@"go/ast".CommentGroup }
	func (@"go/ast".f·2 *@"go/ast".File "esc:0x9") End () (? @"go/token".Pos)
	func (@"go/ast".f·2 *@"go/ast".File "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/ast".f·2.Package }
	type @"go/ast".Package struct { Name string; Scope *@"go/ast".Scope; Imports map[string]*@"go/ast".Object; Files map[string]*@"go/ast".File }
	func (@"go/ast".p·2 *@"go/ast".Package "esc:0x1") End () (? @"go/token".Pos) { return @"go/token".Pos(0x0) }
	func (@"go/ast".p·2 *@"go/ast".Package "esc:0x1") Pos () (? @"go/token".Pos) { return @"go/token".Pos(0x0) }
	func @"".New (@"".pkg·2 *@"go/ast".Package "esc:0xa", @"".importPath·3 string, @"".mode·4 @"".Mode) (? *@"".Package)
	type @"go/ast".Node interface { End() (? @"go/token".Pos); Pos() (? @"go/token".Pos) }
	type @"".Example struct { Name string; Doc string; Code @"go/ast".Node; Play *@"go/ast".File; Comments []*@"go/ast".CommentGroup; Output string; EmptyOutput bool; Order int }
	func @"".Examples (@"".files·2 ...*@"go/ast".File "esc:0x9") (? []*@"".Example)
	func @"".Synopsis (@"".s·2 string "esc:0x1a") (? string)
	var @"".IllegalPrefixes []string
	func @"".init ()
	var @"go/ast".objKindStrings [7]string

$$
_go_.o          0           0     0     644     438782    `
go object linux amd64 go1.6.4 X:none

!
  go13ldio.aregexp.astrings.atext/template.aunicode.aunicode/utf8.ago/ast.ago/token.apath.asort.astrconv.a � "".commentEscape  �
  �
dH�%    H;a��  H��xH��$�   H�D$@    ��$�    tn1�H��H��H9�~aH��$�   H9��J  H��+H��H��H��H��$�   H9��"  H�+�8�u�L$?��`��   ��'��   H��H��H��H9��H�\$@H��H9���   L��$�   H)�H�� tM�H�$    L�D$PL�D$H�l$XH�l$�    H�T$H�L$ H�D$(H��$�   H�$H��$�   H�\$H�T$`H�T$H�L$hH�L$H�D$pH�D$ �    H��x��    H�\$@H��H�D$HH9��8  H9��/  L��$�   H)�H�� tM�H�$    L�D$PL�D$H�l$XH�l$�    H�T$H�L$ H�D$(H��$�   H�$H��$�   H�\$H�T$`H�T$H�L$hH�L$H�D$pH�D$ �    H��$�   H��$�   H��$�   H�D$HH��H�D$@�D$?<'uCH�    H�\$H�    H�\$H�    H�\$H�$H�Z ��H��$�   H�D$HH���B���<`u�H�    H�\$H�    H�\$H�    H�\$H�$H�Z ��H��$�   ��    �    �    �    �U��������$
      �  2runtime.stringtoslicebyte   �  0text/template.HTMLEscape   �  $runtime.panicslice   �  2runtime.stringtoslicebyte   �  0text/template.HTMLEscape   �  "".rdquo   � "".rdquo   �  "".rdquo   �       �	  "".ldquo   �	 "".ldquo   �	  "".ldquo   �
       �
  $runtime.panicslice   �
  $runtime.panicindex   �
  $runtime.panicindex   �
  0runtime.morestack_noctxt   P�  "".autotmp_0014  type.[]uint8 "".autotmp_0013  type.string "".autotmp_0010 /type.[]uint8 "".autotmp_0009 Otype.string "".autotmp_0008  type.int 
"".ch qtype.uint8 "".i _type.int "".last otype.int "".nice @type.bool "".text  type.string "".w  type.io.Writer "������ � f4	
8��66  �� Tgclocals·13bdb4aeeaf63de3cc223d640262ea59 Tgclocals·12fc1489b12fcdedb8fc818b7369b5d9   :$GOROOT/src/go/doc/comment.go�0"".pairedParensPrefixLen  �  �dH�%    H;a��   H��PH�D$`H�D$(    H�D$0H�\$XH�\$@H�D$H1�H�D$8H�\$@H�$H�\$HH�\$H�D$�    H�l$(H�D$�L$ H�� tTH�T$8��(uH�� uH�T$0H��H��H�\$(먃�)u�H��H��H�L$(H�� uH�\$`H�\$0�H�� }�H�T$hH��P�H�\$0H�\$hH��P��    �"�����
      �  &runtime.stringiter2   �  0runtime.morestack_noctxt   0�  "".autotmp_0022  type.int32 "".autotmp_0019 /type.int "".autotmp_0018  type.int "".autotmp_0017  type.int "".autotmp_0016 type.string "".l ?type.int "".parens Otype.int "".~r1  type.int "".s  type.string  ����� � L�	L

%  X� Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·d8fdd2a55187867c76648dc792366181   :$GOROOT/src/go/doc/comment.go�"".emphasize  �  �dH�%    H�D$�H;A��  H��   H��$�   H��$�   H�    H�$H��$�   H�L$H��$�   H�D$�    L��$�   L��$�   H��$�   H��$�   ��$�   H�D$H�L$ H��$�   H�\$(H��$�   H�D$xH�� u$H�<$H�t$L�L$L�D$�T$ �    H�Ĩ   �H�� ��  H�L9���  H�<$H�t$L�L$hL�L$H�\$pH�\$�T$ �    H�T$xH��$�   H�� �q  H�
H��H���Z  H��H�+L��$�   L9��;  H9��2  L��$�   H)�H�� tM�L�D$XL�$H�l$`H�l$�    H�D$H�L$`H9���  H�\$xH��$�    ��  H�H�D$@H��$�   H�H9���  H��$�   H��H�    H�$H�l$hH�l$H�L$pH�L$�    H�\$H�\$xH�\$ H��$�   H�\$(H��$�   H�\$@H�l$`H9��B  H�\$`1�H�D$HH�D$P1ɈL$?H��$�   1�H9�tbH�D$XH�L$`H�    H�$H��$�   H�\$H�D$hH�D$H�L$pH�L$�    H�D$ �\$(H�و\$?H�� ��  H�(H�l$HH�@H�\$xH��$�   ��  H��H�H�� |�� uH�\$XH�\$HH�D$`1ɈL$?H�D$PH�� �]  H�    H�\$H�    H�\$H�    H�\$H��$�   H�$H��$�   H�[ ��H�$    H�\$HH�\$H�\$PH�\$�    H�T$H�L$ H�D$(H��$�   H�$H��$�   H�\$H��$�   H�T$H��$�   H�L$H��$�   H�D$ �    H�    H�\$H�    H�\$H�    H�\$H��$�   H�$H��$�   H�[ ���L$?�� t>H�    H�\$H�    H�\$H�    H�\$H��$�   H�$H��$�   H�[ ��H��$�   H�$H��$�   H�\$H�\$XH�\$H�\$`H�\$��$�   �\$ �    �|$? t>H�    H�\$H�    H�\$H�    H�\$H��$�   H�$H��$�   H�[ ��H�\$PH�� ��   H�    H�\$H�    H�\$H�    H�\$H��$�   H�$H��$�   H�[ ��H�\$xH��$�   v;H��H�H��$�   H9�w L��$�   H)�H�� tM�H��L��������    �    ������    � �:����    �    �    �����    �    �    �    �    �    �N�����������������Z
      d  "".matchRx   �  Pregexp.(*Regexp).FindStringSubmatchIndex   �   "".commentEscape   �   "".commentEscape   �  0"".pairedParensPrefixLen   �  "".matchRx   �  Pregexp.(*Regexp).FindStringSubmatchIndex   �	  ,type.map[string]string   �
  4runtime.mapaccess2_faststr   �  "".html_a   � "".html_a   �  "".html_a   �       �  2runtime.stringtoslicebyte   �  0text/template.HTMLEscape   �  "".html_aq   � "".html_aq   �  "".html_aq   �       �  "".html_i   � "".html_i   �  "".html_i   �       �   "".commentEscape   �  "".html_endi   � "".html_endi   �  "".html_endi   �       �  "".html_enda   � "".html_enda   �  "".html_enda   �       �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `�  &"".autotmp_0034  type.int "".autotmp_0033  type.int "".autotmp_0032 /type.[]uint8 "".autotmp_0031  type.int "".autotmp_0030  type.string "".autotmp_0029  type.string "".autotmp_0028  type.int "".autotmp_0027  type.int "".autotmp_0025  type.int "".autotmp_0024 type.string "".italics �type.bool "".url �type.string "".n �type.int "".match �type.string "".m _type.[]int "".nice Ptype.bool "".words @,type.map[string]string "".line  type.string "".w  type.io.Writer "�����	� � ��/qh]IP+�b!>uC>>>>?ef
 4 T�ur����Fx Tgclocals·2331195bde16ef19bace3004fa98e646 Tgclocals·88f14b8ca07e3b9e0b9cbc5ca8ee0278   :$GOROOT/src/go/doc/comment.go�"".indentLen  �  �dH�%    H;avQH�t$H�L$1�H9�}H9�s4H���� uH��H9�|�H�D$�H9�sH����	u����    �    �    ����������
      �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0   "".~r1  type.int "".s  type.string p p $�! 
 R Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�"".isBlank  �  �dH�%    H;av=H�L$H�� t+H��uH�\$H�� v���
�D$��    �D$ ���D$���    ��������������
      p  $runtime.panicindex   �  0runtime.morestack_noctxt   0   "".autotmp_0039  type.int "".~r1  type.bool "".s  type.string ` ` �8 
 7) Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�"".commonPrefix  �  �dH�%    H;avmL�T$H�|$H�t$ H�T$1�1�H9�}+H9�}&H9�s?H��H9�s,I�,�m @8�uH��H9�|�H9�wH�|$(H�D$0��    �    �    �    �z�������������

      �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `   "".~r2 @type.string "".b  type.string "".a  type.string � � $�%( 
 g) Tgclocals·b4c25e9b09fd0cf9bb429dcefe91c353 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�"".unindent  �  �dH�%    H�D$�H;A�~  H���   H��$�   H�� uH���   �H��$�   H�� �H  H�H�$H�NH�L$�    H�D$H��$�   H��$�    �  L�CL9���  L�I��H�D$xL�D$pH��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$8H��$�   H�l$8H9��  H�t$HH�� ��  H�.H�VH�|$@H��$�   H��$�   H��$�   H�l$PH��$�   H�T$XH�� �E  H���4  H�� �#  �] ��
��< uH�,$H�T$�    H�\$H��$�   H9���  H��$�   H��H�\$pH�$H�\$xH�\$H��$�   H�l$H��$�   H�D$�    H�|$@H�t$HH�\$ H�\$pL�L$(L�L$xH��H��H�l$8H9������L�L$0L��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$8L��$�   H�l$8H9���   L�L$HI�� �  I�1I�QH�L$@H��H�t$`H�T$hH�� ��   H����   H�� ��   ���
��< uvH�\$0H��H��$�   H9���   H)�I��H��$�   H�� tM�H��$�   H��L��L��$�   H��L9�s^H��H�H��$�   H�CH��$�   �=     u H�I��H��H�l$8H9��"���H���   �H�$H�T$�    L�L$HH�L$@���    �    �    1��3���H��   �'���A�������    �    1������H��   �������h����    �    �    �    �`���
      �  "".indentLen   �  "".indentLen   �  "".commonPrefix   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0�  2"".autotmp_0064  type.bool "".autotmp_0063  type.string "".autotmp_0062  type.*string "".autotmp_0061  type.int "".autotmp_0060  type.int "".autotmp_0058 Otype.string "".autotmp_0057 �type.*string "".autotmp_0056 �type.int "".autotmp_0055  type.int "".autotmp_0054  type.string "".autotmp_0053  type.int "".autotmp_0052  type.int "".autotmp_0051  type.[]string "".autotmp_0050  type.string "".autotmp_0049  type.int "".autotmp_0046 /type.[]string "".autotmp_0045  type.int "".autotmp_0044 �type.int "".s �type.string "".s �type.string "".line otype.string "".n �type.int "".line �type.string "".prefix �type.string "".block  type.[]string .��������
 � d�'`pF
c5v

  W�S�w Tgclocals·cb395d89503762333b1bfb09ba74eb12 Tgclocals·6bdcbbfceecc5cba590c8a52e9a888b3   :$GOROOT/src/go/doc/comment.go�"".heading  �	  �	dH�%    H;a�:  H��@1�H�\$XH�\$`H�\$HH�$H�\$PH�\$�    H�T$H�L$H�� u1�H�\$XH�\$`H��@�H�T$HH�$H�L$PH�L$�    �D$�D$,�$�    �\$�� ��  �\$,�$�    �\$�� ��  H�\$HH�$H�\$PH�\$�    �D$�D$,�$�    �\$�� u'�\$,�$�    �\$�� u1�H�\$XH�\$`H��@�H�\$HH�$H�\$PH�\$H�    H�\$H�D$   �    H�\$ H�� |1�H�\$XH�\$`H��@�H�L$HH�D$PH�L$0H�$H�D$8H�D$�D$'   �    H�t$0H�L$8H�D$H�� }H�\$HH�\$XH�\$PH�\$`H��@�H��H��H9�};H��H��H9�syH�.���su$H��H��H9�})H��H��H9�sNH�.��� t1�H�\$XH�\$`H��@�H��H��H��H9�wH)�I��H�� tM�H��L���1����    �    �    1�H�\$XH�\$`H��@��    �������������
      n  "strings.TrimSpace   �  >unicode/utf8.DecodeRuneInString   �   unicode.IsLetter   �  unicode.IsUpper   �  Funicode/utf8.DecodeLastRuneInString   �   unicode.IsLetter   �  unicode.IsDigit   �  Zgo.string.",.;:!?+*/=()[]{}_^°&§~%#@<\">\\"   �   strings.IndexAny   �  "strings.IndexRune   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �	  0runtime.morestack_noctxt   @�  "".autotmp_0073  type.int "".autotmp_0071  type.int "".autotmp_0070  type.int "".autotmp_0069  type.bool "".autotmp_0068  type.bool "".b type.string "".r 'type.int32 "".~r1  type.string "".line  type.string D�D���H�W�V�O � `�#"4
,8
/F%'  6��9 Tgclocals·f47057354ec566066f8688a4970cff5a Tgclocals·d8fdd2a55187867c76648dc792366181   :$GOROOT/src/go/doc/comment.go�"".anchorID  �  �dH�%    H;a��   H��H1�H�\$`H�\$hH�    H�$H�\$PH�\$H�\$XH�\$H�    H�\$H�D$    �    H�L$(H�D$0H�$    H�    H�\$H�D$   H�L$8H�L$H�D$@H�D$ �    H�\$(H�\$`H�\$0H�\$hH��H��    �A����
      L   "".nonAlphaNumRx   �  go.string."_"   �  Bregexp.(*Regexp).ReplaceAllString   �   go.string."hdr-"   �  *runtime.concatstring2   �  0runtime.morestack_noctxt   @�  "".autotmp_0074 type.string "".~r1  type.string "".line  type.string ��� � �#� 
 Wi Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad   :$GOROOT/src/go/doc/comment.go�"".ToHTML  �  �dH�%    H��$(���H;A��  H��X  H��$p  H�$H��$x  H�\$�    H�L$H�D$H�T$ H��$   H��$  H��$  H��$�   H�D$P    H��$�   H�D$HH��$�   H�L$`H�\$PH�l$HH9���  H�\$`H�� �  H�H�sH�SH�kH��$8  H��$@  H��$   H��$H  H��$(  H��$P  H��$0  H��$  H�� ��  H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��H��$   H��$(  H��$0  H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9���   H�D$XH�� ��   H�H�hH�L$@H��$�   H��$�   H��$`  H�$H��$h  H�\$H�T$xH�T$H��$�   H�l$H��$�  H�\$ �D$(�    H�D$XH�L$@H��H��H�l$8H9��o���H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��H�\$`H�� H�\$`H�\$PH��H�\$PH�\$PH�l$HH9�����H��X  É ����H����  H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��1�H��$�   H��$�   H��$   H��$(  H��$0  H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9��t  H�D$XH�� ��  H�H�hH�L$@H��$�   H�T$hH��$�   H�l$pH��$�   H�� ��   H�\$hH�$H�\$pH�\$�    H�L$H�D$H�$    H��$�   H�L$H��$�   H�D$�    H�T$H�L$ H�D$(H��$�   H�T$H��$�   H�L$H��$�   H�D$H��$h  H�$H��$`  H�[ ��H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��H��$`  H�$H��$h  H�\$H�\$hH�\$H�\$pH�\$�D$ �    H�D$XH�L$@H��H��H�l$8H9������H��$�   H�� u>H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ������� ����H������H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ��H��$   H��$(  H��$0  H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9���   H�D$XH�� ��   H�H�hH�L$@H��$�   H��$�   H��$`  H�$H��$h  H�\$H��$�   H�T$H��$�   H�l$H�D$     �D$( �    H�D$XH�L$@H��H��H�l$8H9��p���H�    H�\$H�    H�\$H�    H�\$H��$h  H�$H��$`  H�[ ������� �5����������    �:�������������R
      x  "".blocks   �  "".html_p   � "".html_p   �  "".html_p   �       �  "".emphasize   �  "".html_endp   � "".html_endp   �  "".html_endp   �	       �
  "".html_h   �
 "".html_h   �  "".html_h   �       �  "".anchorID   �  2runtime.stringtoslicebyte   �       �  "".html_hq   � "".html_hq   �  "".html_hq   �       �   "".commentEscape   �  "".html_hq   � "".html_hq   �  "".html_hq   �       �  "".html_endh   � "".html_endh   �  "".html_endh   �       �  "".html_pre   � "".html_pre   �  "".html_pre   �       �  "".emphasize   �  "".html_endpre   � "".html_endpre   �  "".html_endpre   �       �  0runtime.morestack_noctxt   P�  <"".autotmp_0097  type.string "".autotmp_0096  type.*string "".autotmp_0095  type.int "".autotmp_0094  type.int "".autotmp_0093  type.string "".autotmp_0092  type.*string "".autotmp_0091  type.int "".autotmp_0090  type.int "".autotmp_0089 �type.string "".autotmp_0088 �type.*string "".autotmp_0087 �type.int "".autotmp_0086 �type.int "".autotmp_0084 ?type."".block "".autotmp_0083 �type.*"".block "".autotmp_0082 �type.int "".autotmp_0081 �type.int "".autotmp_0080  type.[]string "".autotmp_0079 �type.[]uint8 "".autotmp_0078  type.[]string "".autotmp_0077 �type.[]string "".autotmp_0076 �type.[]"".block "".autotmp_0075 �type.[]"".block "".line �type.string "".line �type.string 
"".id �type.string "".line �type.string "".b type."".block "".words @,type.map[string]string "".text  type.string "".w  type.io.Writer ""������ � ��"�
>sG>.>5
>}"w>7>>+
>sF>721 D ;��`��1�n��`) Tgclocals·46ae46c0833abd65a9bd508c0d4723b4 Tgclocals·a7d2bdfc04e5cad614b789a6f5ec96df   :$GOROOT/src/go/doc/comment.go�"".blocks  �*  �*dH�%    H��$����H;A�M
  H��  1�H��$�  H��$�  H��$�  1�H��$  H��$  H��$   1�H��$�   H��$   H��$  �D$G �D$F 1�H��$X  H��$`  H��$h  H��$X  H�-    H�(H��$�   H�hH��$  H�hH�D$XH��$�  H�$H��$�  H�\$H�    H�\$H�D$   �    H�T$ H�L$(H�D$0H��$(  H�$H��$0  H�L$H��$8  H�D$�    1�H��$0  H9���   H��$(  H��H�t$PL��$0  L9���  H��H�H�3H�SH��$�   H�t$pH��$�   H�T$xH�� ��  H����  H�� ��  ���
��< tjH�T$XH���H�t$PH���D$GH��$0  H9��d���H�T$XH���H��$  H��$�  H��$  H��$�  H��$   H��$�  H�Đ  �H�4$H�T$�    H�t$PH�\$H�� �3  H�T$XH���H�D$PH��$(  H��$0  I��H��H9�}eH��H��H9���  H��H�H�3H��$�   H�KH��$�   H�� ��  H����  H�� ��  ���
���� �*  H��H9�|�L9�~^H��H��H��H9��  H��H�H�3H�t$`H�KH�L$hH�� ��  H����  H�� ��  ���
���� tH��L9��L��$8  L��H��L9���  I9��w  L)�M)�I��I�� tHk�I�H�D$PL��$�   L�$H��$�   H�l$L��$�   L�D$�    H�t$P1�HǄ$p     H��$�   H��$x  H��$�   H��$�  H��$�   H��$�  H��$  H��$  H��$   H��H��H9�wpH��$  H��H��Hk� H�H��$p  H�+H��$�  H�kH��$�  H�kH��$x  �=     uH�k�D$F �����L�CL�$H�l$�    H�t$P��H�-    H�,$H�L$H�D$H�T$H�\$ �    H�t$PH�L$(H�\$0H�T$8H��H��H��$  H��$   H��$  �=����    �    1��G���H��   �;����    H��H��H�D$HH9�sJH��H�H�H�$H�NH�L$�    L�L$PH��$(  H��$0  H�D$HH�\$H�� ������|����    �    1��^���H��   �R����    �|$G �x  �|$F �m  H��$0  H��H��H9��U  H��H��H��$(  L��$0  L9��}  H��H�H�H��$�   H�kH��$�   H�� �I  H���8  H�� �'  ���
��< ��  H��$(  L��$0  H��H��L9���  H��H�H�H��$�   H�kH��$�   H�� ��  H����  H�� ��  ���
��< �|  H��H��$(  H��$0  H��H9��a  H��H�H�H�$H�NH�L$�    H�t$PH�\$H�� �,  H��$�   H�$H��$�   H�\$�    H�t$PH�\$H��$�   H�D$H��$�   H�� ��  H�T$XH���1�H��$x  H��$�  H��$�  HǄ$p     H�    H�$�    H�D$H�� �t  HǄ$H     HǄ$P     H��$@  H��$�   H�hH��$�   �=     �  H�(H��$x  H��$H  H��$�  H��$P  H��$�  H��$  H��$  H��$   H��H��H9�wtH��$  H��H��Hk� H�H��$p  H�+H��$�  H�kH��$�  H�kH��$x  �=     uH�kH�t$PH���D$F�����L�CL�$H�l$�    ��H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$  H��$   H��$  �>���H�$H�l$�    H��$@  ������ �����D$G �D$F H��$(  L��$0  H��L9���   H��H�H�+H��$�   H�kH��$�   H��$�   H��$   H��$  H��H��H9�wRH��$   H��H��Hk�H�H��$�   H�kH��$�   �=     uH�+H������H�$H�l$�    H�t$P��H�-    H�,$H�L$H�D$H�T$H�\$ �    H�t$PH�L$(H�\$0H�T$8H��H��H��$   H��$  H��$�   �[����    ������    �    1��b���H��   �V����    �    1������H��   ������    �    1��^���H��   �R����    �    ������������������Z
      �  "".blocks.func1   �  go.string."\n"   �  $strings.SplitAfter   �  "".unindent   �       �       �  "".indentLen   �	       �  "".unindent   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]"".block   �  "runtime.growslice   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  "".indentLen   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  "".indentLen   �  "".heading   �       �  type.[1]string   �  "runtime.newobject   � (runtime.writeBarrier   �  (runtime.writeBarrier   �!  .runtime.writebarrierptr   �!  type.[]"".block   �"  "runtime.growslice   �#  .runtime.writebarrierptr   �% (runtime.writeBarrier   �&  .runtime.writebarrierptr   �&  type.[]string   �&  "runtime.growslice   �'  $runtime.panicindex   �'  $runtime.panicindex   �(  $runtime.panicindex   �(  $runtime.panicindex   �(  $runtime.panicindex   �)  $runtime.panicindex   �)  $runtime.panicindex   �)  $runtime.panicindex   �)  0runtime.morestack_noctxt   P�  J"".autotmp_0133 �type.string "".autotmp_0131 �type.[]string "".autotmp_0130  type."".block "".autotmp_0128  type.int "".autotmp_0126  type.int "".autotmp_0125 ?type."".block "".autotmp_0123  type.int "".autotmp_0120 ottype.struct { F uintptr; para *[]string; out *[]"".block } "".autotmp_0118  type.int "".autotmp_0116  type.int "".autotmp_0114  type.int "".autotmp_0112  type.int "".autotmp_0111  type.int "".autotmp_0110  type.int "".autotmp_0109  type.int "".autotmp_0108  type.int "".autotmp_0106  type.int "".autotmp_0102  type.int "".autotmp_0101  type.int "".s �type.string "".s �type.string "".s �type.string "".s �type.string "".s �type.string "".head �type.string "".pre �type.[]string "".j �type.int "".line �type.string "".i �type.int "".lines �type.[]string "".close �type.func() """.lastWasHeading �type.bool "".lastWasBlank �type.bool "".para �type.[]string "".out �type.[]"".block "".~r1  type.[]"".block "".text  type.string ""������ � ��<IB+/E
j
8["b[60�98[!�&�G
�	SPx�edbI?% j �:�C!��+<O3�26
3�&@�+<� Tgclocals·3836fb0d9c1e7dd27acd0557fec71b90 Tgclocals·f67a1bd37088b83155134772c74a5fc0   :$GOROOT/src/go/doc/comment.go�"".ToText  �  �dH�%    H��$����H;A�n  H��  1�H��$X  H��$`  ��$h  H��$p  H��$x  H��$�  H��$�  H��$�  H��$�  H��$X  H��$�  H��$`  H��$�  H��$p  H��$�  H��$x  H��$�  H��$�  H��$�  H�$H��$�  H�\$�    H�L$H�D$H�T$ H��$   H��$  H��$  H��$�   H�D$P    H��$�   H�D$HH��$�   H�L$`H�\$PH�l$HH9��A  H�\$`H�� �=  H�H�SH�sH�KH��$8  H��$@  H��$   H��$H  H��$(  H��$P  H��$0  H��$  H�� ��   H��$�   1�H��$�   H�t$8H��$�   H��H�l$8H9�}nH�D$XH�� ��   H�H�hH�L$@H��$�   H��$�   H��$X  H�$H�T$xH�T$H��$�   H�l$�    H�D$XH�L$@H��H��H�l$8H9�|�H��$X  H�$�    H�\$`H�� H�\$`H�\$PH��H�\$PH�\$PH�l$HH9������H�Ę  É �S���H���R  H�    H�\$H�    H�\$H�    H�\$H��$�  H�$H��$�  H�[ ��H��$   H��$(  H��$0  H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9���   H�D$XH�� ��   H�H�hH�L$@H��$�   H��$�   H�$    H��$�   H�T$H��$�   H�l$H�    H�\$H�D$    �    H�\$(H�|$H�H�H�KH�OH��$X  H�$�    H�D$XH�L$@H��H��H�l$8H9��Q���H��$X  H�$�    �n���� �C���H���]���H�    H�\$H�    H�\$H�    H�\$H��$�  H�$H��$�  H�[ ��H��$   H��$(  H��$0  H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9������H�D$XH�� ��  H�H�hH�L$@H��$�   H��$�   H��$�   H�T$hH��$�   H�l$pH�� ��  H����  H�� ��  ���
��< ��   H�$    H�    H�\$H�D$   �    H�T$H�L$ H�D$(H��$�   H�T$H��$�   H�L$H��$�   H�D$H��$�  H�$H��$�  H�[ ��H�D$XH�L$@H��H�������H�$    H��$�  H�\$H��$�  H�\$�    H�T$H�L$ H�D$(H��$�   H�T$H��$�   H�L$H��$�   H�D$H��$�  H�$H��$�  H�[ ��H�$    H��$�   H�\$H��$�   H�\$�    H�T$H�L$ H�D$(H��$�   H�T$H��$�   H�L$H��$�   H�D$H��$�  H�$H��$�  H�[ ��������    1��o���H��   �c���� �����������    �m����������������2
      �  "".blocks   �  ."".(*lineWrapper).write   �	  ."".(*lineWrapper).flush   �
  
"".nl   �
 
"".nl   �
  
"".nl   �       �  go.string."\n"   �  *runtime.concatstring2   �  ."".(*lineWrapper).write   �  ."".(*lineWrapper).flush   �  
"".nl   � 
"".nl   �  
"".nl   �       �  go.string."\n"   �  2runtime.stringtoslicebyte   �       �  2runtime.stringtoslicebyte   �       �  2runtime.stringtoslicebyte   �       �  $runtime.panicindex   �  0runtime.morestack_noctxt   ��  F"".autotmp_0169  type.string "".autotmp_0168  type.*string "".autotmp_0167  type.int "".autotmp_0166  type.int "".autotmp_0165  type.string "".autotmp_0164  type.*string "".autotmp_0163  type.int "".autotmp_0162  type.int "".autotmp_0161 �type.string "".autotmp_0160 �type.*string "".autotmp_0159 �type.int "".autotmp_0158 �type.int "".autotmp_0156 �type."".block "".autotmp_0155 �type.*"".block "".autotmp_0154 �type.int "".autotmp_0153 �type.int "".autotmp_0152  type.[]uint8 "".autotmp_0151  type.[]uint8 "".autotmp_0150 �type.[]uint8 "".autotmp_0147  type.[]string "".autotmp_0146  type.[]string "".autotmp_0145 �type.[]string "".autotmp_0144 �type.[]"".block "".autotmp_0143 �type.[]"".block "".s �type.string "".line �type.string "".line �type.string "".line �type.string "".b �type."".block "".l &type."".lineWrapper "".width �type.int "".preIndent `type.string "".indent @type.string "".text  type.string "".w  type.io.Writer ""������ � ��"�
�
W(.4+
>se
>sIrww	 > ��,��YW��wZ? Tgclocals·a8e198e4544b9f4af27e2179a8f48de0 Tgclocals·da53b597af7c02fca1968f95e2ccd079   :$GOROOT/src/go/doc/comment.go�."".(*lineWrapper).write  �  �dH�%    H�D$�H;A��  H���   H��$�   H�X0H�� uP�X�� tGH�H�hH�    H�\$H�    H�\$H�    H�\$H�l$pH�,$H�L$hH�Y ��H��$�   H��   @�hH��$�   H�$H��$�   H�\$�    H�T$H�D$H�L$ H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$@H��$�   H��H�l$@H9���  H�D$PH�� ��  H�H�hH�L$HH�T$xH��$�   H�T$XH�$H�l$`H�l$�    H��$�   H�L$H�L$8H�X0H�� ~nH�X0H�h8H�H�H�hH9�~WH�H�hH�    H�\$H�    H�\$H�    H�\$H�l$pH�,$H�L$hH�Y ��H��$�   H�@0    H�@8    H�X0H�� ��   H�$    H�X H�|$H�H�H�KH�O�    H�T$H�L$ H�D$(H��$�   H�� ��  H�;H�kH��$�   H�T$H��$�   H�L$H��$�   H�D$H�l$pH�,$H�|$hH�_ ��H��$�   H�X8H�-    H9��%  L�    H��H�8H�hL��$�   L�D$H��$�   H�\$H��$�   H�L$H�l$pH�,$H�|$hH�_ ��H�$    H�\$XH�\$H�\$`H�\$�    H�T$H�L$ H�D$(H��$�   H�� ��   H�;H�kH��$�   H�T$H��$�   H�L$H��$�   H�D$H�l$pH�,$H�|$hH�_ ��H��$�   H�H0H�h8L�D$8L�H�H�h0H�@8   H�D$PH�L$HH��H��H�l$@H9��o���H���   É�i����    ��o���� �Z����    �@���(
      �  
"".nl   � 
"".nl   �  
"".nl   �       �  strings.Fields   �  <unicode/utf8.RuneCountInString   �  
"".nl   � 
"".nl   �  
"".nl   �       �  2runtime.stringtoslicebyte   �	       �	  "".space   �	  "".space   �       �  2runtime.stringtoslicebyte   �       �  $runtime.panicslice   �  0runtime.morestack_noctxt   0�  "".autotmp_0181 �type.string "".autotmp_0180 �type.*string "".autotmp_0179 �type.int "".autotmp_0178 �type.int "".autotmp_0177  type.int "".autotmp_0176  type.[]uint8 "".autotmp_0175  type.[]uint8 "".autotmp_0173 �type.[]uint8 "".autotmp_0172 _type.[]string "".autotmp_0171 /type.[]string "".w �type.int "".f �type.string "".text type.string "".l  (type.*"".lineWrapper  �����
 � f�'G�*!G�`� 
  w��� Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 Tgclocals·77c75893cdd92181c21e4e3e10e9f609   :$GOROOT/src/go/doc/comment.go�."".(*lineWrapper).flush  �  �dH�%    H;avqH��HH�D$PH�X0H�� uH��H�H�H�hH�    H�\$H�    H�\$H�    H�\$H�l$@H�,$H�L$8H�Y ��H�D$PH�@8    H�@0    H��H��    �v���������
      b  
"".nl   z 
"".nl   �  
"".nl   �       �  0runtime.morestack_noctxt   �  "".l  (type.*"".lineWrapper ���X� � $�
D 
 d, Tgclocals·87d20ce1b58390b294df80b886db78bf Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad   :$GOROOT/src/go/doc/comment.go�"".New  �  �dH�%    H��$����H;A��  H��  H��$�   W�H����    H��$�   H�$H��$�  H�\$H��$�  H�\$�    H��$�   H�$�    H��$�   H�$�    H��$0  H�$�    H�\$H��$�   H�\$H��$�   H�\$H��$�   H�    H��   H�    H�$H��$(  H�\$H�L$@H�L$H�D$HH�D$�    H�\$ H�� ��  H�H�KH�kH��$�   H�$H��$�   H�L$H��$�   H�l$�    H�\$H��$�   H�\$ H��$�   H�\$(H��$�   H��$@  H�H�$H�KH�L$H�KH�L$H�D$@   �    H�\$ H��$�   H�\$(H��$�   H�\$0H��$�   H��$X  H�$H��$�  H��H�� �D$�    H�\$H��$�   H�\$H��$�   H�\$ H��$�   H��$@  H�H�$H�KH�L$H�KH�L$H�D$U   �    H�\$ H�\$hH�\$(H�\$pH�\$0H�\$xH��$`  H�$�D$�    H�\$H�\$PH�\$H�\$XH�\$ H�\$`H�    H�$�    H�D$H��$   H�D$8H�� �  H�D$H�\$H�    H�$�    H��$�  H�� ��  H�\$8H�� ��  L�CL�D$H�l$H�-    H�,$�    H�\$8H��$�  H�k(H��$�  �=     �z  H�k H�\$8H��$�   H�k8H��$�   H�k@H��$�   �=     �-  H�k0H��$  H�l$8H�� �
  L�EHL�D$H�\$H�    H�$�    H�\$8H�� ��  H��$(  �=     ��  H�k`H�\$8H��$�   H�kpH��$�   H�kxH��$�   �=     �]  H�khH�\$8H��$�   H���   H��$�   H���   H��$�   �=     �  H���   H�\$8H��$�   H���   H��$�   H���   H��$�   �=     ��   H���   H�\$8H�l$pH���   H�l$xH���   H�l$h�=     ueH���   H�\$8H�l$XH���   H�l$`H���   H�l$P�=     uH���   H�\$8H��$�  H�Ĉ  �L���   L�$H�l$�    ��L���   L�$H�l$�    �L���   L�$H�l$�    �?���L���   L�$H�l$�    �����L�ChL�$H�l$�    ����L�C`L�$H�l$�    �C�����#����E �����L�C0L�$H�l$�    �����L�C L�$H�l$�    �s�����$����E ����� �������&����    �������N
      d�  runtime.duffzero   �  0"".(*reader).readPackage   �  <"".(*reader).computeMethodSets   �  2"".(*reader).cleanupTypes   �  "".sortedKeys   �  go.string."BUG"   �  4type.map[string][]*"".Note   �  4runtime.mapaccess1_faststr   �  "".noteBodies   �  "".sortedValues   �  "".sortedTypes   �  "".sortedValues   �	  "".sortedFuncs   �
  type."".Package   �
  "runtime.newobject   �  type.string   �  (runtime.typedmemmove   �  type.string   �  (runtime.typedmemmove   � (runtime.writeBarrier   � (runtime.writeBarrier   �  type.[]string   �  (runtime.typedmemmove   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   P�  "".autotmp_0196 � type.*"".Package "".autotmp_0195 �type.[]*"".Func "".autotmp_0194 � type.[]*"".Value "".autotmp_0193 �type.[]*"".Type "".autotmp_0192 � type.[]*"".Value "".autotmp_0191 �type.[]string "".autotmp_0190 �type.[]*"".Note "".autotmp_0189 �type.string "".autotmp_0188 �type.[]string "".r �type."".reader "".~r3 @ type.*"".Package "".mode 0type."".Mode "".importPath type.string "".pkg  (type.*go/ast.Package ""��	���� � t�"+
8�VMMI1�5��& N \��MV4.6��
=4 Tgclocals·d40f86804c765b65adbc82845c11e455 Tgclocals·b58df2d7616fbb6904d034404c8af93c   2$GOROOT/src/go/doc/doc.go�"".Examples  �-  �-dH�%    H��$����H;A�+  H��  1�H��$�  H��$�  H��$�  1�H��$  H��$   H��$(  H��$�  H��$�  H��$�  H��$�  1�H��$�  H�D$`H��$�  H��H�l$`H9���  H��$�   H�(H�L$hH�l$x�D$F H�D$H    1�H��$0  H��$8  H��$@  H�\$xH�� �U
  H�KH�C H�k(H��$�  H�D$X    H��$�  H�D$PH��$x  H��$�   H�\$XH�l$PH9���   H��$�   H�� ��	  H�3H�SH��$�   H��$   H��$�   H��H��$�   1�H9�tH�[H�-    H9���	  H��H��   < �  H�YH��K��  H�\$HH��H�\$HH��$�   H��H��$�   H�\$XH��H�\$XH�\$XH�l$PH9��H����|$F ��   H�\$HH����   H��$8  H����   H�\$xH��$�   H�    1�H9��7  H��$�   H��$0  H��$8   �  H�+H�� ��  H��$�   H�E H��$�   �=     ��  H�M(H�\$xH�$�    H�D$H��$0  H��$8   ��  H�+H�� �z  �=     �V  H�E0H��$  H��$   H��$(  H��H��$P  H��$8  H�H)�H�� ~KH�    H�$H��$H  H�t$H�T$H��$X  H�D$H�L$ �    H�t$(H�\$0H��$P  H�D$8H�    H�$H��$   H��$   L��$8  L�I��H��$X  H9���  H9���  H)�I)�I��H��$H  I�� tM��H�l$L�D$L�L$H��$0  H�\$ H��$8  H�\$(H��$@  H�\$0�    H��$X  H��$   H��$8  H�H9��  H��H��$H  H��$  H��$   H��$(  H��$�   H�L$hH��H��H�l$`H9��G���H��$  H��$`  H��$   H��$h  H��$(  H��$p  H�    H�$H�    H�\$H�    H�\$H��$`  H�\$H�D$     �    H�\$(H�H�$H�KH�L$�    H��$  H��$�  H��$   H��$�  H��$(  H��$�  H�Ĩ  ��    �    L�E0L�$H�D$�    �����E �~����    L�E(L�$H�L$�    �)����E ������    H�    H�$H�    H�\$H�    H�\$�    H�D$����H��1�H9�tH�[H�-    H9��e  H��H��   < �����H�\$HH��H�\$HH��$�   H�iH�� �(  H�MH�EH��$�   H�$H��$�   H�D$H�    H�\$H�D$   �    �\$ �� ��  H��$�   H�$H��$�   H�\$H�    H�\$H�D$	   �    �\$ �� ��  H��$�   H�$H��$�   H�\$H�    H�\$H�D$   �    H��$�   �\$ �� u�����1�H��$�   H��$�   H�1�H9�t.H�)H�,$�    H��$�   H�\$H��$�   H�\$H��$�   H�i H�,$H�t$xH�� ��  H�^hH�|$H�H�H�KH�OH�KH�O�    H�\$ H��$�   H�\$(H��$�   �\$0�\$GH��$�   H����  H��$�   H��H�� tH��H��$  H��$  H�\$xH�$H��$�   H�k H�l$�    H�\$H��$�   H��$8  H�\$pH�    H�$�    H�\$H��$�   H��$�   H��$  H�kH��$  �=     ��  H�+H��$�   H��$�   H�kH��$�   �=     ��  H�kH�    1�H9��?  H��$�   H�K H��$�   H�� �  H��$�   H�C H��$�   �=     ��  H�K(H��$�   H�� ��  H��$�   �=     ��  H�k0H�\$xH�� �  H�khH��$�   H�� �b  L�C8L�D$H�l$H�-    H�,$�    H��$�   H��$�   H�hXH��$�   �=     ��   H�hPH��H�� ��   L��$�   I�� ��   �l$G@�k`H�l$pH�hhH��$�   H��$0  H��$8  H��$@  H��H��H9�w8H��$8  H��H��$�   �=     uH�+�����H�$H�l$�    �����H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�D$0H�T$8H��H��H��$8  H��$@  H��$0  �z���1��3���� ����L�@PL�$H�l$�    H��$�   ������������z���L�C0L�$H�l$�    �T�����4���L�C(L�$H�L$�    ����������H�    H�$H�    H�\$H�    H�\$�    H�D$����L�CL�$H�l$�    �f���H�$H�l$�    �&����    ������D$F�����E �����1�1�����1�1��`�����
���������    ����x
      �  (type.*go/ast.GenDecl   �  @go.itab.*go/ast.File.go/ast.Node   �	 (runtime.writeBarrier   �
  $"".playExampleFile   � (runtime.writeBarrier   �  $type.[]*"".Example   �  &runtime.growslice_n   �   type.*"".Example   �  ,runtime.typedslicecopy   �  *type."".exampleByName   �  &type.sort.Interface   �  Ngo.itab."".exampleByName.sort.Interface   �  runtime.convT2I   �  sort.Sort   �  $runtime.panicslice   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  "type.*go/ast.File   �   type.go/ast.Node   �  @go.itab.*go/ast.File.go/ast.Node   �   runtime.typ2Itab   �  *type.*go/ast.FuncDecl   �   go.string."Test"   �  "".isTest   �  *go.string."Benchmark"   �  "".isTest   �  &go.string."Example"   �  "".isTest   �  6go/ast.(*CommentGroup).Text   �   "".exampleOutput   �  "".playExample   �  type."".Example   �  "runtime.newobject   �  (runtime.writeBarrier   �! (runtime.writeBarrier   �!  Jgo.itab.*go/ast.BlockStmt.go/ast.Node   �" (runtime.writeBarrier   �# (runtime.writeBarrier   �$  6type.[]*go/ast.CommentGroup   �$  (runtime.typedmemmove   �$ (runtime.writeBarrier   �& (runtime.writeBarrier   �'  .runtime.writebarrierptr   �'  $type.[]*"".Example   �'  "runtime.growslice   �)  .runtime.writebarrierptr   �)  .runtime.writebarrierptr   �*  .runtime.writebarrierptr   �*  ,type.*go/ast.BlockStmt   �*   type.go/ast.Node   �+  Jgo.itab.*go/ast.BlockStmt.go/ast.Node   �+   runtime.typ2Itab   �+  .runtime.writebarrierptr   �+  .runtime.writebarrierptr   �,  $runtime.panicslice   �-  0runtime.morestack_noctxt   `�  L"".autotmp_0226  type.int "".autotmp_0225 �$type.[]*"".Example "".autotmp_0224  type.*uint8 "".autotmp_0222 � type.*"".Example "".autotmp_0221   type.*"".Example "".autotmp_0220 � type.go/ast.Decl "".autotmp_0219 �"type.*go/ast.Decl "".autotmp_0218 �type.int "".autotmp_0217 �type.int "".autotmp_0216 �"type.*go/ast.File "".autotmp_0215 �$type.**go/ast.File "".autotmp_0214 �type.int "".autotmp_0213 �type.int "".autotmp_0212 �*type."".exampleByName "".autotmp_0211  "type.*go/ast.File "".autotmp_0210  "type.*go/ast.File "".autotmp_0209  type.int "".autotmp_0208  type.int "".autotmp_0207  "type.*go/ast.File "".autotmp_0206 �type.string "".autotmp_0205  type.bool "".autotmp_0202  type.int "".autotmp_0200 �type.int "".autotmp_0198 _$type.[]go/ast.Decl "".autotmp_0197 /&type.[]*go/ast.File "".hasOutput �type.bool "".output �type.string "".doc �type.string "".name �type.string "".f �*type.*go/ast.FuncDecl "".decl � type.go/ast.Decl "".flist �$type.[]*"".Example "".numDecl �type.int "".hasTests �type.bool "".file �"type.*go/ast.File "".list �$type.[]*"".Example "".~r1 0$type.[]*"".Example "".files  &type.[]*go/ast.File ""��	����
 � �^<]	�F4D,pH�Y"^�8AA(�E$
.^8,�	�p1K?@?@VW
	
			
 h ���W*��z*��)RK4/
	J Tgclocals·a0565663444d773a05e50b742a3936f2 Tgclocals·57f34913b4e4f52cd021da0277a0692e   :$GOROOT/src/go/doc/example.go� "".exampleOutput  �  �dH�%    H;a��  H��X1�1�H��$�   H��$�   H�\$`H�$H�\$hH�\$H�\$pH�\$H�\$xH�\$�    H�D$(1�H9��7  H�$�    H�L$H�D$H�    H�$H�L$0H�L$H�D$8H�D$�    H�D$H�L$ H�\$(H�\$PH�� ��   H��H�D$@H��H�L$H��   H��H�H�l$8H9���   L�D$0H)�H�� tM�L�D$0L�$H�l$8H�l$H�    H�\$H�D$   �    H�L$ H�D$(H�� ~PH�� vL���
uBH��H��r2H��H��H�� tH��H��H��H��$�   H��$�   Ƅ$�   H��X��    ���    �    �    1�H��$�   H��$�   Ƅ$�    H��X��    �9������������
      �  "".lastComment   �  6go/ast.(*CommentGroup).Text   �  "".outputPrefix   �  @regexp.(*Regexp).FindStringIndex   �  go.string." "   �   strings.TrimLeft   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   p�  "".autotmp_0235  type.int "".loc /type.[]int "".text Otype.string 
"".ok `type.bool "".output @type.string "".comments 6type.[]*go/ast.CommentGroup "".b  ,type.*go/ast.BlockStmt  ����<� � @�+<B>7  RG�� Tgclocals·5cbd57cf8f9b35eac9551b20a42afe1f Tgclocals·fad3647538fe088c3f63d28bb4a0e2d7   :$GOROOT/src/go/doc/example.go�"".isTest  �  �dH�%    H;a�  H��XL�L$hH�|$xL�T$`L�T$(L�D$pL�D$8L�L$0H�|$@I9���   L9���   H9���   L�T$HL�$H�|$PH�|$L�D$H�|$�    L�L$hH�|$x�\$ H��< uƄ$�    H��X�I9�uƄ$�   H��X�L��L9�wNL�D$`H)�H�� tM�8L�D$HL�$H�l$PH�l$�    �\$�$�    �\$H��H����$�   H��X��    1��y����    1��k����    ��������
      �   runtime.eqstring   �  >unicode/utf8.DecodeRuneInString   �  unicode.IsLower   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   P�  "".autotmp_0244  type.bool "".autotmp_0243  type.string "".autotmp_0242  type.int "".autotmp_0241  type.int "".autotmp_0240  type.int "".autotmp_0239 type.string "strings.prefix·3 ?type.string strings.s·2 _type.string "".~r2 @type.bool "".prefix  type.string "".name  type.string 8������U��� � ,�!q6   w� Tgclocals·1c5a071f4ad97fe89533b360c694a573 Tgclocals·709a14768fab2805a378215c02f0d27f   :$GOROOT/src/go/doc/example.go�("".exampleByName.Len      H�\$H�\$ ������ @   "".~r0 0type.int "".s  *type."".exampleByName   �  Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/example.go�*"".exampleByName.Swap  �  �dH�%    H;a��   H��H�T$8H�L$ H�D$(H9���   H��H�+H�l$H9�s~H��L�D$@I9�siJ�,�L�E �=     u>L�H�l$@H9�s*H��H�l$�=     uH�+H���H�$H�l$�    ���    H�$L�D$�    H�L$ H�D$(��    �    �    �    �*�������������
      � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   P0  "".autotmp_0247  type.*"".Example "".j @type.int "".i 0type.int "".s  *type."".exampleByName 0n/0F/ � 
��  �) Tgclocals·3260b5c802f633fd6252c227878dd72a Tgclocals·0c8aa8e80191a30eac23f1a218103f16   :$GOROOT/src/go/doc/example.go�*"".exampleByName.Less  �  �dH�%    H;av{H��(H�T$0H�D$8H�l$HH9�s\H�4�H�.H�M H�$H�MH�L$H�l$PH9�s3H�4�H�.H�|$H�M H�H�MH�O�    H�\$ H�� �D$XH��(��    �    �    �l���������������

      �  "runtime.cmpstring   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `P  "".~r2 Ptype.bool "".j @type.int "".i 0type.int "".s  *type."".exampleByName PhOPO � 
�� 
 d< Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/example.go�"".playExample  �~  �~dH�%    H��$����H;A�{  H��  H��$�  H�kH�� �V  H�}H��$`  H�MH�5    H��$p  H��   H��$h  H��$x  H9��  H��H)�H��H9���  H)�I��H�� tM�H9���  L��$�  L�$H��$�  H�l$H�t$H�D$�    �\$ H��< uHǄ$�      H�Ę  �H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H��$�  H�� �>  H�KH�C H�k(H��$�  1�H��$�  H�D$pH��$�  H��H�l$pH9��  H��$@  H�� ��  H�H�hH�T$xH��$0  H��$8  H��$`  H�$H��$h  H�l$�    H��$`  H��$h  �L$���~���  H��1�H9�tH�[H�-    H9��h  H��H��   �� ��  �D$GH�    H�$H��$�   H�\$H�hH�l$H�|$ �u  H�D$H�\$GH�\$�    H��$@  H�T$xH��H��H�l$pH9������H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H�    H�$�    H�D$H��$P  �  H�    H�$�    H�\$H��$X  H�    H�$�    H�D$H�-    H�(H��$   H��$X  �=     �n  H�hH�� �Y  H��$�   �=     �%  H�hH�� �  H��$�   �=     ��  H�hH�� ��  H��$P  �=     ��  H�h H��$X  �=     �g  H�H��$�  H��$H  H�    1�H9��  H��$H  H��$@  H�$H��$H  H�L$H��$X  H�+H�l$�    H��$P  ��� tHǄ$�      H�Ę  �H��$�   H��$(  W�H����    H�    H�$H�D$H��$(  H�\$�    H��$(  1�H9��E  H��$(  H�� �L  H�H�kH��$   H��$  H�    H�$H�    H�\$H��$�  H�L$H��$�  H�l$�    H�\$ �+@�� ��  H��$   H��$  H�    H�$H�    H�\$H��$�  H�L$H��$�  H�D$�    H�\$ �+@�� �F  H��$   H��$  H�    H�$H�    H�\$H��$�  H�L$H��$�  H�D$�    H�\$ �+@�� ��  H��$(  H�$�    H��$(  1�H9������1�H��$�  ��$�  ��$�  ��$�  H��$�  H��$�  H��$�  H��$�  H��$�  W�H����    H�    H�$H�D$    H��$�  H�\$H��$�  H�\$�    H�\$ H��$�   1�H��$�  H��$�  H��$�  H��$�  H�� �  H�S8H�C@H�kHH��$H  1�H��$@  H�D$pH��$8  H��H�l$pH9���   H��$  H�(H�L$xH��$�   H�]H�� ��  H�kH�M H�$H�MH�L$�    H�T$H��$�  H�L$H��$�  H�D$ H�\$(H��$(  H��$   H�� ��  H��$  H�L$xH��H��H�l$pH9��`���H��$�   1�H9�tH�H�� ~HǄ$�      H�Ę  �E1�L��$�  M��L��$�  M��L��$�  H��$�  H��$�  H��$�  H��$x  E1�H��$p  H�D$xH��$h  H�l$xI9���   H��$8  H�� ��  H�/H�GL�d$pH��$P  H��$X  H��$�  H��$�  E1�L9�tH�mL�    L9���  H�0H��$�   1�H9�t4L��L��L��H��L9���  I��H��$�  H���=     ��  H�3H��I��H�l$xI9��K���H��$�  H�� �v  H�{hH�CpH�kxH��$0  E1�H��$(  H�D$xH��$   H�l$xI9��  H��$  H�7L�d$pH��$�  H�H�� �  H�H�FH�nH��$   H��$�  H�� H��$�  ��  H�*H�m H9���   H��$�   H�NH��H�H�FH�nH��$   H��$�  H��$�  H9���  H��H�H�HH�H�H��H��$�  H�C H��H9�4L��L��L��H��L9���  I��H��$�  H���=     ��  H�3H��I��H�l$xI9������H��$�  H�$L�\$L�T$L�L$�    H�\$ H��$�  H�\$(H��$�  H�\$0H��$�  H�\$8H��$�  H�    H�$�    H�D$1�H�(H�hH�hH�hH�h H�h(H�h0H�h8H�@K   H�@   H�@8   H��$�   H��$�   H��$�  W�H����    H�    H�$H�D$H��$�  H�\$�    H��$�  1�H9��w  H��$�  H�� �_  H�H�SH��$�  H�� �?  H�+H��$  H�kH��$  H��$�  H��$�  H��$�  H�$H��$�  H�T$�    H�\$H��$�  H�\$H��$�  H�    H�$�    H�D$H��$  1�H�(H�hH�hH�hH�h H�    H�$�    H�D$1�H�(H�hH�hH�hH��$�   H��$�  H�hH��$�  �=     �@
  H�hH��$  H�� �#
  �=     ��	  H�CH��$  H��$�   H��$�  H�$H��$�  H�\$�    H��$  H�T$H�D$H9���  H��$�  H�$H��$�  H�D$H��$  H�l$H�L$�    H��$  �\$ �� ��  H��$�   H��$  H�    1�H9��^  H��$  H��$X  H��$P  H��$�   H�S H�k(H�K0H��H��H9���  H�k(H��H��Hk�H�H��$P  H�+H��$X  �=     �E  H�kH��$�  H�$�    H��$�  1�H9������H��$�   H�� �  H�s H�{(H�C0H��$h  H��$p  H��$x  H��H��$  H��$�  H�H)�H�� ~SH�    H�$H��$  H�t$H�|$H��$  H�D$H�L$ �    H��$p  H�t$(H�\$0H��$  H�D$8H�    H�$L��$�  H��H��L�I��H��$  H9��7  H9��.  H)�I)�I��H��$  I�� tHk�I�H�l$L�D$L�L$H��$�  H�\$ H��$�  H�\$(H��$�  H�\$0�    H��$  H��$p  H��$�  H�H9���  H��H��$�   H�C(H�K0H��$  �=     �k  H�k H�    H��$�  HǄ$�     H�    H�$�    H�D$H�     H��$(  H��$�  H�hH��$�  �=     ��  H�h1�H�hH��$�   H�    H�$�    H�D$1�H�(H�hH�hH�hH�h H��$�   H��$�   �=     �x  H�hH�    H�$�    H�D$H��$�   1�H�(H�hH�hH�    H�$�    H�D$1�H�(H�hH�hH�hH�h H��$�   H�� �  �=     ��  H�CH��$�   H�� ��  H��$�   �=     ��  H�kH��$�   H�� �}  H��$�  �=     �Q  H�k H��$�   H��$�   H�    H��$�  HǄ$�     H�    H�$�    H�D$H�     H��$(  H��$�  H�hH��$�  �=     ��  H�h1�H�hH��$�   H��$�   H��$   H��$�   H��$�   H�    H�$�    H�|$H��H�� �c  W��    H��$�   H�� �B  H��$�   �=     �  H�hH�    H�$�    H�\$H�� ��  HǄ$�     HǄ$�     H��$�  H�    1�H9���  H��$   H��$�  H��$`  H�H��$h  �=     �A  H�KH�    1�H9���   H��$�   H��$�  H��H��$`  H�H��$h  �=     ��   H�KH��$�   H��$�  H�k H��$�  H�k(H��$�  �=     ueH�kH��$�   H��$�  H�kpH��$�  H�kxH��$�  �=     uH�khH��$�   H��$�  H�Ę  �L�ChL�$H�l$�    ��L�CL�$H�l$�    �L�CL�$H�L$�    �?���H�    H�$H�    H�\$H�    H�\$�    H�D$�����L�CL�$H�L$�    ����H�    H�$H�    H�\$H�    H�\$�    H�D$�F��������L�@L�$H�l$�    ������ ���������L�@L�$H�l$�    H��$(  �'���L�C L�$H�l$�    ������|���L�CL�$H�l$�    �S�����3���L�CL�$H�D$�    �
���������L�@L�$H�l$�    �u���L�@L�$H�l$�    H��$(  �����L�C L�$H�l$�    �����    �    ������L�CL�$H�l$�    ����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H��$�   H�� tQH��H�l$HH��H�k(H�K0H��$�   �=     u	H�S �	���L�C L�$H�T$�    H��$�   H�D$H�������H�    H�$H�    H�\$H�    H�\$�    H�D$�p���H��$  H��$�  H��$�  H�    H�$�    H�D$H�     H��$(  H��$�  H�hH��$�  �=     uEH�h1�H�hH��$�   H�� t)�=     u	H�C�����L�CL�$H�D$�    �������L�@L�$H�l$�    H��$(  �L�CL�$H�D$�    �����������L�@L�$H�l$�    H��$�   ��������������H�$H�t$�    L�d$pL��$�  L��$�  L��$�  H��$  �@���H�-    H�,$H�L$H�D$L�L$H�\$ �    L�d$pH��$  H��$�   L�\$(L�T$0L�L$8L��I��L��$�  L��$�  L��L��$�  �����    �    �����������H�$H�t$�    L�d$pH��$8  L��$�  L��$�  L��$�  �$���H�-    H�,$H�L$H�D$L�L$H�\$ �    L�d$pH��$8  H��$�   L�\$(L�T$0L�L$8L��I��L��$�  L��$�  L��L��$�  ����H�,$L�D$L�    L�L$�    �����H�$H�L$�    H��$�   H�\$H��$�  H�\$H��$�  H�X1�H9��  H�hH�� �,  H�]H��$�  H�]H��$�  H��$�  H��$�  H��$�  H��uYH�$H��$�  H�D$H�-    H�l$H�D$   �    H��$�  H��$�  �\$ �� tHǄ$�      H�Ę  �H��$�  H���g  H�$H�D$H�-    H�l$H�D$   �    �\$ �� �6  H��$�   H��$  H�    1�H9���   H��$  H��$X  H��$P  H��$�  H��$�  H��$�  H��H��H9�wQH��$�  H��H��Hk�H�H��$P  H�+H��$X  �=     u	H�k����L�CL�$H�l$�    �q���H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�\$0H�T$8H��H��H��$�  H��$�  H��$�  �a���H�    H�$H�    H�\$H�    H�\$�    H�D$�����H��$�  H��$�  H�    H�$H��$�   H�\$H��$�  H�D$H��$�  H�L$�    H�\$ �+@�� ��   H��$�  H��$�  H��$�  H��$�  H��$�  H��$p  H��$�  H��$x  H�    H�$H��$�   H�\$H��$�  H�\$H��$p  H�\$�    H��$�  H��$�  H��$�  H��$�  H�    H�$H��$�   H�\$H��$�  H�\$�    �����������E �������^���������H��$   H��$�  H��$  H��$�  H�    H�$H��$�   H�\$H��$�  H�\$�    ����������H�    H�$H�    H�\$H�    H�\$�    H�D$����H�$H�D$�    ����L�@ L�$H�l$�    H��$   �R���� �2���L�@L�$H�l$�    H��$   �	���� �����L�@L�$H�l$�    H��$   ������ ����L�@L�$H�l$�    H��$   �w����%    ��������f[�����H��1�H9�tH�[H�-    H9��o  H��H��   �� �W���H��H�� �H  H�H H�@(H�k0H��$x  1�H��$p  H�D$XH��$h  H��H�l$XH9�����H��$8  H�� ��  H�H�hH�T$`H��$�  H��$�  H��$P  H�$H��$X  H�l$�    H��$P  H��$X  �T$��Z�v3�  H��1�H9�tH�[H�-    H9��r  H��H��   < ��   H�� ��   H�QH�AH�iH��$`  1�H��$X  H�D$PH��$P  H��H�l$PH9�}mH��$0  H�(H�L$h�D$GH�    H�$H��$�   H�\$H�l$H�|$ tLH�D$H�\$GH�\$�    H��$0  H�L$hH��H��H�l$PH9�|�H��$8  H�T$`H��H�������%    뫉�2���������u�H��1�H9�tH�[H�-    H9�u`H��H��   �� t��D$GH�    H�$H��$�   H�\$H�hH�l$H�|$ tH�D$H�\$GH�\$�    �^����%    ��1�1��1�1������ ����� ����1�1�����1�1������ ���������1��R����    1��D����E �����    �`����
      �  "go.string."_test"   �   runtime.eqstring   �  8type.map[*go/ast.Object]bool   �  runtime.makemap   �  $runtime.ifacethash   �  *type.*go/ast.FuncDecl   �  8type.map[*go/ast.Object]bool   �	  $runtime.mapassign1   �	  (type.map[string]bool   �
  runtime.makemap   �
  type.bool   �
  "runtime.newobject   �  6type.func(go/ast.Node) bool   �  "runtime.newobject   �  �type.struct { F uintptr; inspectFunc *func(go/ast.Node) bool; unresolved map[string]bool; topDecls map[*go/ast.Object]bool; usesTopDecl *bool }   �  "runtime.newobject   �  ("".playExample.func1   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  Jgo.itab.*go/ast.BlockStmt.go/ast.Node   �  go/ast.Inspect   ��  runtime.duffzero   �  (type.map[string]bool   �  &runtime.mapiterinit   �  (type.map[string]bool   �  &"".predeclaredTypes   �  4runtime.mapaccess1_faststr   �  (type.map[string]bool   �  ."".predeclaredConstants   �  4runtime.mapaccess1_faststr   �  (type.map[string]bool   �  &"".predeclaredFuncs   �  4runtime.mapaccess1_faststr   �  &runtime.mapiternext   ��  runtime.duffzero   �  ,type.map[string]string   �  runtime.makemap   �  strconv.Unquote   �   .type.*go/ast.ImportSpec   �! (runtime.writeBarrier   �' (runtime.writeBarrier   �(  *"".stripOutputComment   �)  &type.go/ast.GenDecl   �)  "runtime.newobject   �*�  runtime.duffzero   �+  ,type.map[string]string   �+  &runtime.mapiterinit   �-  strconv.Quote   �.  ,type.go/ast.ImportSpec   �.  "runtime.newobject   �.  (type.go/ast.BasicLit   �.  "runtime.newobject   �/ (runtime.writeBarrier   �0 (runtime.writeBarrier   �1  path.Base   �2   runtime.eqstring   �3  Lgo.itab.*go/ast.ImportSpec.go/ast.Spec   �4 (runtime.writeBarrier   �5  &runtime.mapiternext   �7  $type.[]go/ast.Spec   �7  &runtime.growslice_n   �8   type.go/ast.Spec   �:  ,runtime.typedslicecopy   �; (runtime.writeBarrier   �;   go.string."main"   �<  "type.go/ast.Ident   �<  "runtime.newobject   �= (runtime.writeBarrier   �=  (type.go/ast.FuncDecl   �=  "runtime.newobject   �> (runtime.writeBarrier   �>  (type.go/ast.FuncType   �?  "runtime.newobject   �?  *type.go/ast.FieldList   �?  "runtime.newobject   �@ (runtime.writeBarrier   �A (runtime.writeBarrier   �A (runtime.writeBarrier   �B   go.string."main"   �B  "type.go/ast.Ident   �B  "runtime.newobject   �C (runtime.writeBarrier   �D   type.go/ast.File   �D  "runtime.newobject   �E�  runtime.duffzero   �E (runtime.writeBarrier   �E  &type.[2]go/ast.Decl   �F  "runtime.newobject   �F  Fgo.itab.*go/ast.GenDecl.go/ast.Decl   �G (runtime.writeBarrier   �H  Hgo.itab.*go/ast.FuncDecl.go/ast.Decl   �H (runtime.writeBarrier   �I (runtime.writeBarrier   �J (runtime.writeBarrier   �K  .runtime.writebarrierptr   �K  .runtime.writebarrierptr   �K  .runtime.writebarrierptr   �L  *type.*go/ast.FuncDecl   �L   type.go/ast.Decl   �L  Hgo.itab.*go/ast.FuncDecl.go/ast.Decl   �L   runtime.typ2Itab   �M  .runtime.writebarrierptr   �M  (type.*go/ast.GenDecl   �M   type.go/ast.Decl   �M  Fgo.itab.*go/ast.GenDecl.go/ast.Decl   �M   runtime.typ2Itab   �N  .runtime.writebarrierptr   �N  .runtime.writebarrierptr   �O  .runtime.writebarrierptr   �O  .runtime.writebarrierptr   �P  .runtime.writebarrierptr   �P  .runtime.writebarrierptr   �Q  .runtime.writebarrierptr   �Q  .runtime.writebarrierptr   �Q  $runtime.panicslice   �Q  $runtime.panicslice   �R  .runtime.writebarrierptr   �R  $type.[]go/ast.Spec   �S  "runtime.growslice   �S (runtime.writeBarrier   �T  .runtime.writebarrierptr   �T  .type.*go/ast.ImportSpec   �U   type.go/ast.Spec   �U  Lgo.itab.*go/ast.ImportSpec.go/ast.Spec   �U   runtime.typ2Itab   �V  "type.go/ast.Ident   �V  "runtime.newobject   �V (runtime.writeBarrier   �W (runtime.writeBarrier   �W  .runtime.writebarrierptr   �X  .runtime.writebarrierptr   �X  .runtime.writebarrierptr   �Y  .runtime.writebarrierptr   �Y  .runtime.writebarrierptr   �Z  6type.[]*go/ast.CommentGroup   �[  "runtime.growslice   �\  $runtime.panicindex   �\  $runtime.panicindex   �\  .runtime.writebarrierptr   �]  6type.[]*go/ast.CommentGroup   �^  "runtime.growslice   �_   type.go/ast.Spec   �_  (runtime.panicdottype   �`  path.Base   �b  go.string."."   �b   runtime.eqstring   �c  go.string."_"   �d   runtime.eqstring   �d  Lgo.itab.*go/ast.ImportSpec.go/ast.Spec   �f (runtime.writeBarrier   �f  .runtime.writebarrierptr   �g  $type.[]go/ast.Spec   �g  "runtime.growslice   �h  .type.*go/ast.ImportSpec   �h   type.go/ast.Spec   �h  Lgo.itab.*go/ast.ImportSpec.go/ast.Spec   �i   runtime.typ2Itab   �i  (type.map[string]bool   �j  4runtime.mapaccess1_faststr   �k  ,type.map[string]string   �l  $runtime.mapassign1   �m  (type.map[string]bool   �m  "runtime.mapdelete   �n  (type.map[string]bool   �o  "runtime.mapdelete   �o  ,type.*go/ast.BlockStmt   �o   type.go/ast.Node   �o  Jgo.itab.*go/ast.BlockStmt.go/ast.Node   �p   runtime.typ2Itab   �p  .runtime.writebarrierptr   �p  .runtime.writebarrierptr   �q  .runtime.writebarrierptr   �q  .runtime.writebarrierptr   �r  .runtime.writebarrierptr   �s  (type.*go/ast.GenDecl   �v  $runtime.ifacethash   �w  ,type.*go/ast.ValueSpec   �x  8type.map[*go/ast.Object]bool   �y  $runtime.mapassign1   �{  *type.*go/ast.TypeSpec   �{  8type.map[*go/ast.Object]bool   �|  $runtime.mapassign1   �~  $runtime.panicslice   �~  0runtime.morestack_noctxt   0�  �"".autotmp_0353  type.*uint8 "".autotmp_0352  type.*uint8 "".autotmp_0350  $type.[]go/ast.Decl "".autotmp_0349 �"type.*go/ast.File "".autotmp_0348  $type.*go/ast.Ident "".autotmp_0347  $type.*go/ast.Ident "".autotmp_0345 �*type.*go/ast.FuncType "".autotmp_0344 �*type.*go/ast.FuncDecl "".autotmp_0343  $type.*go/ast.Ident "".autotmp_0342  $type.*go/ast.Ident "".autotmp_0341  type.int "".autotmp_0340 �
$type.[]go/ast.Spec "".autotmp_0339  $type.[]go/ast.Spec "".autotmp_0338  type.*uint8 "".autotmp_0337   type.go/ast.Spec "".autotmp_0336  $type.*go/ast.Ident "".autotmp_0335  $type.*go/ast.Ident "".autotmp_0334 �*type.*go/ast.BasicLit "".autotmp_0333  .type.*go/ast.ImportSpec "".autotmp_0332  type.string "".autotmp_0331 �(type.*go/ast.GenDecl "".autotmp_0330  "type.go/token.Pos "".autotmp_0329  "type.go/token.Pos "".autotmp_0328  "type.go/token.Pos "".autotmp_0325 �4type.**go/ast.CommentGroup "".autotmp_0324  type.int "".autotmp_0323  type.int "".autotmp_0322   type.go/ast.Spec "".autotmp_0321  "type.*go/ast.Spec "".autotmp_0320  type.int "".autotmp_0319  type.int "".autotmp_0318  type.*uint8 "".autotmp_0317   type.go/ast.Spec "".autotmp_0316  type.string "".autotmp_0315 �.type.*go/ast.ImportSpec "".autotmp_0314 �0type.**go/ast.ImportSpec "".autotmp_0313  type.int "".autotmp_0312  type.int "".autotmp_0311 �:type.map.bucket[string]string "".autotmp_0310 �4type.map.hdr[string]string "".autotmp_0308 ��type.*struct { F uintptr; inspectFunc *func(go/ast.Node) bool; unresolved map[string]bool; topDecls map[*go/ast.Object]bool; usesTopDecl *bool } "".autotmp_0307 �$type.*go/ast.Ident "".autotmp_0306 �&type.**go/ast.Ident "".autotmp_0305 �type.int "".autotmp_0304  type.int "".autotmp_0303  type.uint32 "".autotmp_0301   type.go/ast.Spec "".autotmp_0300 � type.go/ast.Spec "".autotmp_0299 �"type.*go/ast.Spec "".autotmp_0298  type.int "".autotmp_0297  type.int "".autotmp_0295  type.bool "".autotmp_0294   type.go/ast.Decl "".autotmp_0293 � type.go/ast.Decl "".autotmp_0292 �"type.*go/ast.Decl "".autotmp_0291  type.int "".autotmp_0290  type.int "".autotmp_0288  *type.*go/ast.FuncDecl "".autotmp_0287  (type.*go/ast.GenDecl "".autotmp_0286  .type.*go/ast.ImportSpec "".autotmp_0285  type.string "".autotmp_0284  type.string "".autotmp_0283 �6type.map.iter[string]string "".autotmp_0281  type.int "".autotmp_0280  type.int "".autotmp_0279 �	6type.[]*go/ast.CommentGroup "".autotmp_0278  $type.[]go/ast.Spec "".autotmp_0277  type.int "".autotmp_0276  type.string "".autotmp_0275 �type.string "".autotmp_0274  type.string "".autotmp_0273  type.bool "".autotmp_0272  type.string "".autotmp_0271  .type.*go/ast.ImportSpec "".autotmp_0270 �	2type.[]*go/ast.ImportSpec "".autotmp_0269 �type.string "".autotmp_0267 �type.string "".autotmp_0266  type.bool "".autotmp_0265 �type.string "".autotmp_0264  type.bool "".autotmp_0263  type.string "".autotmp_0262 �2type.map.iter[string]bool "".autotmp_0260 �,type.*go/ast.BlockStmt "".autotmp_0259  type.bool "".autotmp_0258 �	(type.[]*go/ast.Ident "".autotmp_0257  type.bool "".autotmp_0256 �$type.[]go/ast.Spec "".autotmp_0255 �type.bool "".autotmp_0254 �$type.[]go/ast.Decl "".autotmp_0253 �type.string "".autotmp_0252 �type.int "".autotmp_0251 �type.int "".autotmp_0250 �type.int "".autotmp_0249 �type.int "".autotmp_0248 �type.int "".&usesTopDecl �type.*bool "".&inspectFunc �8type.*func(go/ast.Node) bool "".~r0 �$type.*go/ast.Ident go/ast.name·2 �type.string "".~r0 �$type.*go/ast.Ident go/ast.name·2 �type.string go/ast.name·2 �type.string "strings.suffix·3 �type.string strings.s·2 �type.string "".funcDecl �*type.*go/ast.FuncDecl "".s �.type.*go/ast.ImportSpec "".p �type.string "".n �type.string "".importDecl �(type.*go/ast.GenDecl "".c �2type.*go/ast.CommentGroup "".c �2type.*go/ast.CommentGroup "".s � type.go/ast.Spec "".comments �6type.[]*go/ast.CommentGroup "".n �type.string "".err �type.error "".p �type.string "".s �.type.*go/ast.ImportSpec "".blankImports �
$type.[]go/ast.Spec "".namedImports �,type.map[string]string "".n �type.string "".unresolved �(type.map[string]bool "".spec � type.go/ast.Spec "".decl � type.go/ast.Decl "".topDecls �8type.map[*go/ast.Object]bool "".~r2  "type.*go/ast.File "".body ,type.*go/ast.BlockStmt "".file  "type.*go/ast.File Z"������������������
 �? ��"�8lG"&8 �.Xj�$�^\"2!|64\�4T>
���	$�0J:I*!�0<:; *+��8GCHQ	
�-Z6YZ]=3n	3n30&K	C��YwJ%
J2/.-r%=g~R?		1C	
 � ���M �
br����D��*2����{WK*�wU�
-I#%<
'"
)\>2m)NO%Nd�c�)ZQ�Jj4L���W	  Tgclocals·ab21a96c86932eb21e674bd4000cfd30 Tgclocals·0b5e8d15b1b34de9bb59946bbdd0aacd   :$GOROOT/src/go/doc/example.go�$"".playExampleFile  �  �dH�%    H��$H���H;A�9  H��8  H��$@  H�� �  H�ShH��$  H�KpH�kxH��$  H��$  H�� ��   H�� ��  H�*H�,$�    L�D$H�t$L��$�   H�=    H��$�   H��	   H��$�   H��$�   H9���  H9��v  H9��f  L��$�   L�$H��$�   H�D$H�|$H�D$�    �\$ H��< tJH��$  H��$  H���  H��H��L��$  H�� tI��H��$  H��$  L��$  1�H��$�   H��$�   H��$   H��$@  H�� ��  H�KH�C H�k(H��$0  H�D$H    H��$(  H�D$@H��$   H�L$`H�\$HH�l$@H9���  H�\$`H�� �N  H�H�kH��$�   H��$�   H��$�   H��$�   H��$�   1�H9�tH�[H�-    H9���  H��$�   H��   < ��  H�L$PH�YH�� ��  H�kH�M H�$H�MH�L$H�    H�\$H�D$   �    �\$ �� ��  H�    H�$�    H�D$H�\$PH�� �]  H�D$pH�D$H�\$H�    H�$�    H�    H��$�   HǄ$�      H�    H�$�    H�D$H�     H�D$XH��$�   H�hH��$�   �=     ��  H�h1�H�hH�\$p�=     ��  H�CH�\$PH�k H�,$H��$  H�\$H��$  H�\$H��$  H�\$�    H�D$ H�\$(H��$  H�\$0H��$  H�\$8H��$  H�\$p�=     �   H�C H�\$pH�\$hH�    1�H9���  H�\$hH��$�   H��$�   H��$�   H��$�   H��$   H��H��H9��  H��$�   H��H��Hk�H�H��$�   H�+H��$�   �=     ��  H�kH�\$`H��H�\$`H�\$HH��H�\$HH�\$HH�l$@H9��F���H�    H�$�    H�D$H��$@  H�� �p  H�D$xH�D$H�\$H�    H�$�    H�    H��$�   HǄ$�      H�    H�$�    H�D$H�     H�D$XH��$�   H�hH��$�   �=     ��   H�h1�H�hH�\$x�=     ��   H�CH�\$xH��$�   H�k H��$   H�k(H��$�   �=     u_H�kH�\$xH��$  H�kpH��$  H�kxH��$  �=     uH�khH�\$xH��$H  H��8  �L�ChL�$H�l$�    ��L�CL�$H�l$�    �L�CL�$H�D$�    �H���L�@L�$H�l$�    H�D$X���������L�CL�$H�l$�    ����H�-    H�,$H�L$H�D$H�T$H�\$ �    H�L$(H�D$0H�T$8H��H��H��$�   H��$   H��$�   ����H�    H�$H�    H�\$H�    H�\$�    H�D$� ���L�C L�$H�D$�    �����L�CL�$H�D$�    �[���L�@L�$H�l$�    H�D$X�#���������������/���1�1������������K����    1�������    1������    �������    ������b
      �  6go/ast.(*CommentGroup).Text   �  *go.string."Copyright"   �   runtime.eqstring   �  *type.*go/ast.FuncDecl   �	  &go.string."Example"   �	  "".isTest   �
  (type.go/ast.FuncDecl   �
  "runtime.newobject   �
  (type.go/ast.FuncDecl   �
  (runtime.typedmemmove   �   go.string."main"   �  "type.go/ast.Ident   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   �  *"".stripOutputComment   � (runtime.writeBarrier   �  Hgo.itab.*go/ast.FuncDecl.go/ast.Decl   � (runtime.writeBarrier   �   type.go/ast.File   �  "runtime.newobject   �   type.go/ast.File   �  (runtime.typedmemmove   �   go.string."main"   �  "type.go/ast.Ident   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $type.[]go/ast.Decl   �  "runtime.growslice   �  *type.*go/ast.FuncDecl   �   type.go/ast.Decl   �  Hgo.itab.*go/ast.FuncDecl.go/ast.Decl   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt    �  8"".autotmp_0397  $type.*go/ast.Ident "".autotmp_0396  $type.*go/ast.Ident "".autotmp_0393 �$type.*go/ast.Ident "".autotmp_0392  $type.*go/ast.Ident "".autotmp_0391 � type.go/ast.Decl "".autotmp_0390 �"type.*go/ast.Decl "".autotmp_0389  type.int "".autotmp_0388  type.int "".autotmp_0386  *type.*go/ast.FuncDecl "".autotmp_0385  type.bool "".autotmp_0384 �*type.*go/ast.FuncDecl "".autotmp_0383 /$type.[]go/ast.Decl "".autotmp_0382  type.string "".autotmp_0379 �type.int "".autotmp_0378 �type.string "".autotmp_0377 �type.int 
"".&f �"type.*go/ast.File "".&newF �*type.*go/ast.FuncDecl go/ast.name·2 �type.string go/ast.name·2 �type.string "strings.prefix·3 �type.string strings.s·2 �type.string "".f �*type.*go/ast.FuncDecl "".d � type.go/ast.Decl "".decls �$type.[]go/ast.Decl "".comments _6type.[]*go/ast.CommentGroup "".~r1 "type.*go/ast.File "".file  "type.*go/ast.File ""������ � ��".�J��C07{1`.F}22V2
	 ^ s�3+��
6+�#)Z96 Tgclocals·93d42c534c9b7817c9d67e4a28433e4e Tgclocals·6cf11449797bbc22c96eb58e2aa7d4d6   :$GOROOT/src/go/doc/example.go�*"".stripOutputComment  �  �dH�%    H�D$�H;A��  H���   1�H��$  H��$  H��$  H��$�   H�$H��$�   H�\$H��$�   H�\$H��$�   H�\$�    H�\$ H�\$HH�D$(1�H9���  H�D$XH�$�    H�L$H�D$H�    H�$H�L$hH�L$H�D$pH�D$�    �\$�� ��  H�\$XH�� ��  H�H�CH�kH��$�   H��$�   H�� H��$�   �R  H�)H�m H�l$@H�    H�$�    H��$�   H�D$H�� �  H�)H�(H�iH�D$`L�@L�D$H�l$H�-    H�,$�    H�D$`H�l$@H�h H�D$PH��$�   H��H�    H�$H�D$H�D$�    L�L$H�|$ H�t$(H�\$HH��$�   H9���  L��$�   H��H�    H�$L�L$xL�L$H��$�   H�|$H��$�   H�t$L��$�   L�D$ H��$�   H�T$(H��$�   H�l$0�    H�D$HH��$�   L��$�   H9���   L�L$xH)�I)�I�� tM��I��L��L��H��H��H��$�   L��$�   H9���   L��$�   H)�I)�I�� tM��H�    H�$H��$�   H�t$L��$�   L�T$H��$�   H�|$L��$�   L�L$ H��$�   H�l$(L��$�   L�D$0�    H�\$PH��$   H�\$xH��$  H��$�   H��$  H��$�   H��$  H���   ��    �    �    � ������    ��s���H��$�   H��$   H��$�   H��$  H��$�   H��$  H��$�   H��$  H���   ��    �=����������������(
      �  "".lastComment   �  6go/ast.(*CommentGroup).Text   �  "".outputPrefix   �  8regexp.(*Regexp).MatchString   �  *type.go/ast.BlockStmt   �  "runtime.newobject   �  $type.[]go/ast.Stmt   �  (runtime.typedmemmove   �  6type.[]*go/ast.CommentGroup   �  "runtime.makeslice   �  2type.*go/ast.CommentGroup   �  ,runtime.typedslicecopy   �
  2type.*go/ast.CommentGroup   �  ,runtime.typedslicecopy   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   ��  "".autotmp_0410 �,type.*go/ast.BlockStmt "".autotmp_0408 _6type.[]*go/ast.CommentGroup "".autotmp_0407  type.int "".autotmp_0406  6type.[]*go/ast.CommentGroup "".autotmp_0405 /6type.[]*go/ast.CommentGroup "".autotmp_0402 �type.string "".~r0 �"type.go/token.Pos "".newComments �6type.[]*go/ast.CommentGroup "".newBody �,type.*go/ast.BlockStmt "".last �2type.*go/ast.CommentGroup "".i �type.int "".~r3 P6type.[]*go/ast.CommentGroup "".~r2 @,type.*go/ast.BlockStmt "".comments 6type.[]*go/ast.CommentGroup "".body  ,type.*go/ast.BlockStmt  ����q� � P�9GUe,	
4��B	H * l(�D8��� Tgclocals·87c30dc0786889497a80d853dd7fef3f Tgclocals·0ce45eb4af445847db003d38f23f3ab0   :$GOROOT/src/go/doc/example.go�"".lastComment  �  �dH�%    H;a��   H�T$H�D$0    H�D$(    L�"L�Z I��H�T$L�T$H�\$ 1�L9�}2H�
H�� tqH�9H�qH�iH�� vYH�/H�] L9�}H��H��L9�|��H�yH��H�H�qH�iH9�s"H��H�3H�~H�H�L9��H�D$(H�L$0��    �    ���    �.�����������������
      �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `   "".autotmp_0425  "type.go/token.Pos "".autotmp_0424  "type.go/token.Pos "".autotmp_0423  "type.go/token.Pos "".autotmp_0417  "type.go/token.Pos "".autotmp_0415  type.int "".last P2type.*go/ast.CommentGroup "".i @type.int "".c 6type.[]*go/ast.CommentGroup "".b  ,type.*go/ast.BlockStmt � � 4�*
#	-
  �* Tgclocals·d98f60bd8519d0c68364b2a1d83af357 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/example.go�$"".filterIdentList  �  �dH�%    H;a�E  H��X1�H�\$xH��$�   H��$�   1�H�t$H�T$`H�D$hH�\$pH�\$P1�H�D$HH�D$ H�T$@H��H�l$ H9���   H�D$8H�(H�L$(H�l$0H�� ��   H�]H�H�$H�KH�L$�    H�t$�\$�� ��   H�\$`L�D$hL9���   H��H�l$0�=     uZH�+H��H�t$H�D$8H�L$(H��H��H�l$ H9��i���H�l$pH9�wL�D$`L�D$xH��$�   H��$�   H��X��    H�$H�l$�    H�t$��    듉E �/����    ������������������
      �  "go/ast.IsExported   � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `�  "".autotmp_0435 ?&type.**go/ast.Ident "".autotmp_0434 otype.int "".autotmp_0433 _type.int "".autotmp_0432  (type.[]*go/ast.Ident "".autotmp_0429 /(type.[]*go/ast.Ident "".x O$type.*go/ast.Ident "".j type.int "".~r1 0(type.[]*go/ast.Ident "".list  (type.[]*go/ast.Ident  ����-� � :$.C;(0  ��) Tgclocals·adb3347b296419e60da36d67f8b7ce43 Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0   :$GOROOT/src/go/doc/exports.go�$"".hasExportedName  �  �dH�%    H;a��   H��@H�T$HH�D$PH�\$XH�\$81�H�D$0H�D$H�T$(H��H�l$H9�}EH�D$ H�(H�L$H�,$�    �\$�� t
�D$`H��@�H�D$ H�L$H��H��H�l$H9�|��D$` H��@��    �^�����������������
      �  4go/ast.(*Ident).IsExported   �  0runtime.morestack_noctxt   @�  "".autotmp_0441 ?&type.**go/ast.Ident "".autotmp_0440 _type.int "".autotmp_0439 Otype.int "".autotmp_0437 /(type.[]*go/ast.Ident "".~r1 0type.bool "".list  (type.[]*go/ast.Ident �[�$ � >?


 
 ZV Tgclocals·f47057354ec566066f8688a4970cff5a Tgclocals·83ead081cd909acab0dcd88a450c1878   :$GOROOT/src/go/doc/exports.go�&"".removeErrorField  �
  �
dH�%    H�D$�H;A�O  H��   H��$�   H�kH�� �*  H�]H�\$hH�]H�\$pH�]H�\$xH�D$0    H�L$hH�D$pH�\$xH��$�   H�D$@    H��$�   H�D$8H��$�   H�L$PH�\$@H�l$8H9���   H�\$PH��D$/H�jH�� utH�T$HH�Z H�H�$H�KH�L$�    H�T$HH�L$H�L$XH�D$H�D$`H��u7H�$H�D$H�-    H�l$H�D$   �    H�T$H�\$ �� t�D$/ �|$/ t9H�\$hH�l$0L�D$pL9��  H��=     ��   H�H�\$0H��H�\$0H�\$PH��H�\$PH�\$@H��H�\$@H�\$@H�l$8H9�����H�D$pH�\$0H9�}H��$�   H��   @�kH�\$0H�l$xH9�wnL�D$hH��H��$�   H��H�kH�� tLH��$�   H�MH��$�   H�EL��L��$�   �=     uH�]H�Ę   �L�EL�$H�\$�    ��E ��    H�$H�T$�    �����    �E ������    �������������������
      �  "".baseTypeName   �  "go.string."error"   �   runtime.eqstring   � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicslice   �	  .runtime.writebarrierptr   �	  $runtime.panicindex   �	  0runtime.morestack_noctxt   �  "".autotmp_0449 �&type.**go/ast.Field "".autotmp_0448 �type.int "".autotmp_0447 �type.int "".autotmp_0446  (type.[]*go/ast.Field "".autotmp_0445  type.int "".autotmp_0443 /(type.[]*go/ast.Field "".fname type.string "".keepField �type.bool "".field �$type.*go/ast.Field "".j �type.int "".list _(type.[]*go/ast.Field "".ityp  4type.*go/ast.InterfaceType  ����B� � bX1	U
o,.\  ��
( Tgclocals·37a2283f5c69c342946cad8073b58fca Tgclocals·82a1413d9c726b969ce192c6dcea957e   :$GOROOT/src/go/doc/exports.go�8"".(*reader).filterFieldList  �  �dH�%    H�D$�H;A�  H���   Ƅ$   H��$  1�H9�uH���   �H��$  H�� ��  H�kH��$�   H�kH��$�   H�kH��$�   H�D$P    H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$`H��$�   H��H�l$`H9��_  H��$�   H� H�L$h�D$G H�hH�l$HH�� �V  H��$�   H�$H��$   H�\$H��$�   H�X H�|$H�H�H�KH�O�    H�L$ H�D$(H��$�   H�$H��$�   H�D$�    H��$�   �\$�� �y  �D$G�|$G ��   H��$�   H�$H�D$    H��$�   H�� �;  H�^ H�|$H�H�H�KH�O�    H��$�   H�l$PL��$�   L9���   H��H��$�   �=     ��   H�+H�\$PH��H�\$PH��$�   H�L$hH��H��H�l$`H9������H��$�   H�\$PH9�}Ƅ$  H�\$PH��$�   H9�wiL��$�   H��H��$  H�� tLH��$�   H�KH��$�   H�kL��L��$�   �=     uH�kH���   �L�CL�$H�l$�    ����    H�$H�l$�    �"����    �����H��$  1�H9��y���H���o���H��$�   H�,$H�L$H�-    H�l$H�D$   �    �\$ �� �6����D$GH��$�   H��$  H�\$pH��H�D$xH�PxH���   H���   H��H��H9�w4H���   H��H�l$p�=     uH�+�����H�$H�l$�    �����H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H�\$xH�� tWH��H�l$XH��H���   H���   H��$�   �=     u	H�Sx�b���L�CxL�$H�T$�    H��$�   H�D$X�>�����H��$�   H�XH�H�$H�KH�L$H�KH�L$�    H�T$H�L$ H�D$(H��$�   H�� ��   H��$�   H�KH��$�   H�CH��$�   �=     uEH�SH��$�   H�[H�l$HH9�})Ƅ$  H��$�   H�kH�� ~
�D$G�x����s�����L�CL�$H�T$�    뫉�w�����2����    �������������,
      �  B"".(*reader).recordAnonymousField   �  "go/ast.IsExported   �  ."".(*reader).filterType   � (runtime.writeBarrier   �
 (runtime.writeBarrier   �
  .runtime.writebarrierptr   �
  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  "go.string."error"   �   runtime.eqstring   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  8type.[]*go/ast.InterfaceType   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $"".filterIdentList   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   P�  ,"".autotmp_0461 �&type.**go/ast.Field "".autotmp_0460 �type.int "".autotmp_0459 �type.int "".autotmp_0458  (type.[]*go/ast.Field "".autotmp_0457  type.int "".autotmp_0456  type.int "".autotmp_0455  type.int "".autotmp_0453 _(type.[]*go/ast.Ident "".autotmp_0451 /(type.[]*go/ast.Field "".typ �4type.*go/ast.InterfaceType "".r �type.*"".reader "".fname �type.string "".n �type.int "".keepField �type.bool "".field �$type.*go/ast.Field "".j �type.int "".list �(type.[]*go/ast.Field  "".removedFields @type.bool "".ityp 04type.*go/ast.InterfaceType "".fields  ,type.*go/ast.FieldList "".parent $type.*"".namedType "".r  type.*"".reader .�������� �
 ��'6	XG4"C:3":[!VV�x
! 6 �(i�

	Q�_@� Tgclocals·ba362c851cf6718bcf08a64a3f3a3743 Tgclocals·b6cb89307147056cbbf19b02d7f6310a   :$GOROOT/src/go/doc/exports.go�8"".(*reader).filterParamList  �  �dH�%    H;a��   H��PH�D$`1�H9���   H��H�� ��   H�PH�@H�kH�l$H1�H�D$@H�D$ H�T$8H��H�l$ H9�}\H�D$0H�(H�L$(H�\$XH�$H�D$    H�� t<H�] H�|$H�H�H�KH�O�    H�D$0H�L$(H��H��H�l$ H9�|�H��PÉE 뿉 �d����    �&���������
      �  ."".(*reader).filterType   �  0runtime.morestack_noctxt    �  "".autotmp_0469 ?&type.**go/ast.Field "".autotmp_0468 _type.int "".autotmp_0467 Otype.int "".autotmp_0466 /(type.[]*go/ast.Field "".fields ,type.*go/ast.FieldList "".r  type.*"".reader  ����� � (�I4  �A Tgclocals·2f2d69f12d345ece4be5273d9b84f0bb Tgclocals·83ead081cd909acab0dcd88a450c1878   :$GOROOT/src/go/doc/exports.go�."".(*reader).filterType  �  �dH�%    H;a�,  H��XH�L$pH�D$xH�L$HH�$H�D$PH�D$�    H�|$hH�t$`H�T$HH�L$P�D$=Bj	���  =�Z�Q��   =Ns;/u/H��1�H9�tH�[H�-    H9���   H��   �� tH��X�=�Z�Qu�H��1�H9�tH�[H�-    H9���   H��   < t�H�4$H�D$    H�L$8H�� t^H�YH�|$H�H�H�KH�O�    H�\$`H�$H�D$    H�t$8H�� t!H�^H�|$H�H�H�KH�O�    �Y�����ۉ�1�1��y���1��<���=;�5�ufH��1�H9�tH�[H�-    H9���   H��H��   �� t9H�4$H�D$    H�� t!H�]H�|$H�H�H�KH�O�    ������E ��=Bj	������H��1�H9�tH�[H�-    H9�uXH��   < �����H�4$H�|$H�L$@H�iH�l$H�D$    �    �\$ �� tH�\$@H��   @�k�\����W���1�1��1�1��6���==�O���   =���ufH��1�H9�tH�[H�-    H9���   H��H��   �� t9H�4$H�D$    H�� t!H�]H�|$H�H�H�KH�O�    ������E ��==�O������H��1�H9�tH�[H�-    H9�uXH��H��   �� �����H�4$H�|$H�hH�l$H�D$0H�D$�    �\$ �� tH�\$0H��   @�k�X����S���1�1��1�1��6���=���ueH��1�H9�tH�[H�-    H9���   H��H��   �� t8H�4$H�l$(H�mH�l$�    H�\$`H�$H�\$(H�kH�l$�    �����=�z�������H��1�H9�tH�[H�-    H9�uKH��H��   �� �����H�4$H�D$    H�� t!H�XH�|$H�H�H�KH�O�    �l���� ��1�1��1�1��D����    �����������(
      j  $runtime.ifacethash   �  $type.*go/ast.Ident   �  (type.*go/ast.MapType   �  ."".(*reader).filterType   �  ."".(*reader).filterType   �  ,type.*go/ast.ParenExpr   �  ."".(*reader).filterType   �  .type.*go/ast.StructType   �  8"".(*reader).filterFieldList   �	  ,type.*go/ast.ArrayType   �
  ."".(*reader).filterType   �  4type.*go/ast.InterfaceType   �  8"".(*reader).filterFieldList   �  *type.*go/ast.FuncType   �  8"".(*reader).filterParamList   �  8"".(*reader).filterParamList   �  *type.*go/ast.ChanType   �  ."".(*reader).filterType   �  0runtime.morestack_noctxt   @�  "".autotmp_0473  type.go/ast.Expr "".autotmp_0472  type.bool "".autotmp_0471  type.bool "".t ?(type.*go/ast.MapType "".t O4type.*go/ast.InterfaceType "".t _*type.*go/ast.FuncType "".t /.type.*go/ast.StructType "".typ   type.go/ast.Expr "".parent $type.*"".namedType "".r  type.*"".reader "������ � ���0/0&49%D/('4/
/N/$#8+
/C/8,/+ . 4�9��c~	� Tgclocals·948a0e540dd9ee4dc893ee9411d99e55 Tgclocals·54334d948b35c5006059bc936ec0efb4   :$GOROOT/src/go/doc/exports.go�."".(*reader).filterSpec  �  �dH�%    H�D$�H;A�1  H���   H��$�   H��$�   H��$�   H�$H��$�   H�D$�    H��$�   H��$�   �D$=�u:H��1�H9�tH�[H�-    H9���  H��   �� tƄ$  H���   �=Z�v3�/  H��1�H9�tH�[H�-    H9��n  H��H��   �� ��   H�T$8H�� ��   H�ZH�H�$H�KH�L$H�KH�L$�    H�|$8H�T$H�L$ H�D$(H�� ��   H��$�   H�OH��$�   H�GH��$�   �=     u_H�WH�oH�� ~AH��$�   H�$H�D$    H�_ H�|$H�H�H�KH�O�    Ƅ$  H���   �Ƅ$   H���   �L�GL�$H�T$�    H�|$8댉�X��������=����u�H��1�H9�tH�[H�-    H9��/  H��H��   < t�H�L$@H�iH�� �  H�MH�EH�L$xH�$H��$�   H�D$�    H��$�   �\$�� �u  H��$�   H�\$HH�\$@H�kH�� �M  H�MH��$�   H�EH��$�   H�� tGH����   H�$H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� tN1�H��$�   H�$H�D$H�t$@H�� t,H�^H�|$H�H�H�KH�O�    Ƅ$  H���   É��H�    H�$H�\$HH�k`H�l$H��$�   H�L$H��$�   H�D$�    H�D$ �\$(H�(�� tH���b���H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$pH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$hH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$`H�    H�$�    H�|$H��H�� ��  W�H����    H�D$PH��$�   H�hH��$�   �=     �2  H�hH�� �  H�l$p�=     ��   H�h0H�� ��   H�l$h�=     ��   H�hPH�� ��   H�l$`�=     umH�hXH��$�   H��$�   H��$�   H��$�   H�D$0H�D$XH�    H�$H�\$HH�k`H�l$H��$�   H�\$H�\$XH�\$�    H�D$0����L�@XL�$H�l$�    H�D$P�{���� �b���L�@PL�$H�l$�    H�D$P�<���� ����L�@0L�$H�l$�    H�D$P������ �����L�@L�$H�l$�    H�D$P������y����E ����H�������H�l$xH�,$H�L$H�-    H�l$H�D$   �    �\$ �� �����H��$�   H��   @�kp�}����E �����1�1������1�1�����1��D����    �����������������J
      �  $runtime.ifacethash   �  .type.*go/ast.ImportSpec   �  ,type.*go/ast.ValueSpec   �  $"".filterIdentList   � (runtime.writeBarrier   �  ."".(*reader).filterType   �  .runtime.writebarrierptr   �  *type.*go/ast.TypeSpec   �	  "go/ast.IsExported   �
  go.string."_"   �   runtime.eqstring   �  ."".(*reader).filterType   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".namedType   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  "go.string."error"   �   runtime.eqstring   �  0runtime.morestack_noctxt   P�  ("".autotmp_0489 �$type.*"".namedType "".autotmp_0485 � type.go/ast.Spec "".autotmp_0484 �$type.*"".namedType "".autotmp_0483 otype.string "".autotmp_0482 �"type."".methodSet "".autotmp_0481 �"type."".methodSet "".autotmp_0480 �&type."".embeddedSet "".autotmp_0479 Otype.string "".autotmp_0478  type.bool "".autotmp_0476 /(type.[]*go/ast.Ident "".typ �$type.*"".namedType "".name �type.string "".r �type.*"".reader "".name �type.string "".s �*type.*go/ast.TypeSpec "".s �,type.*go/ast.ValueSpec "".~r2 @type.bool "".tok 0&type.go/token.Token "".spec  type.go/ast.Spec "".r  type.*"".reader J�������������� � d�s<
|
1	3L��@ R H��2~�TLz5�
###Kc Tgclocals·d696fea639189e6f0ee17af9ebd01687 Tgclocals·cb1549917f9fe0533af2fa9f39272c98   :$GOROOT/src/go/doc/exports.go� "".copyConstType  �  �dH�%    H;a�V  H��h1�H��$�   H��$�   H�L$pH�D$xH�L$XH�$H�D$`H�D$�    H�t$XH�T$`�L$��Ns;/�  H��1�H9�tH�[H�-    H9���  H�T$(H��   < ��   H�    H�$�    H�D$1�H�(H�hH�hH�hH�\$(H�� ��   H�kH�D$@L�@L�D$H�l$H�-    H�,$�    H�D$@H��$�   H�(H�D$@H�    1�H9�tH�\$@H��$�   H��$�   H��h�H�    H�$H�    H�\$H�    H�\$�    H�D$뷉�f������+�e��  H��1�H9�tH�[H�-    H9���  H��H��   �� ��  H��H�(E1�L9�tH�mL�    L9���  H�SH��   H�T$0�� �R  H�hH�� �<  H�]H�\$HH�]H�\$PH�    H�$�    H�D$H�     H�D$@H�l$PH�hH�l$H�=     ��  H�h1�H�hH�D$ H�    H�$�    H�D$1�H�(H�hH�hH�hH�\$0H�� ��  H�kH�D$@L�@L�D$H�l$H�-    H�,$�    H�D$@H��$�   H�(H�D$@H�    H�$�    H�\$H�\$8H�\$8H�� �  H�l$ �=     ��   H�kH�    1�H9���   H�L$@H�\$8H�� ��   H�D$XH�H�L$`�=     ueH�KH�\$8H�\$8H�    1�H9�tH�\$8H��$�   H��$�   H��h�H�    H�$H�    H�\$H�    H�\$�    H�D$�L�CL�$H�L$�    닉�j���H�    H�$H�    H�\$H�    H�\$�    H�D$�$���L�CL�$H�l$�    �������������r���L�@L�$H�l$�    H�D$@�����E ����1�H��$�   H��$�   H��h�1�1�����1�1��A���H�D$(    1��&����    �����������������N
      �  $runtime.ifacethash   �  $type.*go/ast.Ident   �  "type.go/ast.Ident   �  "runtime.newobject   �  type.string   �  (runtime.typedmemmove   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �  $type.*go/ast.Ident   �   type.go/ast.Expr   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �   runtime.typ2Itab   �  2type.*go/ast.SelectorExpr   �  $type.*go/ast.Ident   �  "type.go/ast.Ident   �  "runtime.newobject   � (runtime.writeBarrier   �	  "type.go/ast.Ident   �	  "runtime.newobject   �
  type.string   �
  (runtime.typedmemmove   �
  0type.go/ast.SelectorExpr   �  "runtime.newobject   � (runtime.writeBarrier   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   � (runtime.writeBarrier   �  Pgo.itab.*go/ast.SelectorExpr.go/ast.Expr   �  2type.*go/ast.SelectorExpr   �   type.go/ast.Expr   �  Pgo.itab.*go/ast.SelectorExpr.go/ast.Expr   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  $type.*go/ast.Ident   �   type.go/ast.Expr   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   P�  &"".autotmp_0504  type.*uint8 "".autotmp_0503  type.*uint8 "".autotmp_0502 _2type.*go/ast.SelectorExpr "".autotmp_0501  $type.*go/ast.Ident "".autotmp_0500  $type.*go/ast.Ident "".autotmp_0499  $type.*go/ast.Ident "".autotmp_0497 O$type.*go/ast.Ident "".autotmp_0494  type.go/ast.Expr "".autotmp_0493  2type.*go/ast.SelectorExpr "".autotmp_0492  $type.*go/ast.Ident "".autotmp_0491  $type.*go/ast.Ident "".autotmp_0490  $type.*go/ast.Ident "".~r0 �$type.*go/ast.Ident go/ast.name·2 ?type.string 
"".id o$type.*go/ast.Ident "".typ $type.*go/ast.Ident "".~r2 0 type.go/ast.Expr "".pos  "type.go/token.Pos "".typ   type.go/ast.Expr <����������"� �1�X t�)n�=;5�1��%X-M��
	 . F\L�KL�JAg Tgclocals·0f0d539f72a0076bd99eb5022e35364d Tgclocals·e4ca007442f0c3cdda096ebe56a943a8   :$GOROOT/src/go/doc/exports.go:$GOROOT/src/go/doc/example.go�6"".(*reader).filterSpecList  �  �dH�%    H�D$�H;A�  H���   1�H��$   H��$  H��$  H��$�   H��@��  1�H�|$pH��H�|$xH��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$0H��$�   H��H�l$0H9��p  H�D$HH�� �c  H�H�@H�T$8H��$�   H��$�   H�D$XH�\$P1�H9�tH�[H�-    H9��  H��H�h H�� ��   H�� ��   H�T$@H��H�� ��  H�RH�CH�kH��$�   H��$�   H�� H��$�   ��  H�*H�m H�$H�|$H�l$�    H�T$@H�L$H�D$ H�� �c  H��$�   H�J H��$�   �=     �&  H�B(H�T$@H�� �  H�ZH�H�$H�KH�L$H�KH�L$�    �\$�� ��  1�H�|$pH��H�|$xH�D$HH�T$8H��H��H�l$0H9������1�H�T$(H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$0H��$�   H��H�l$0H9���   H�D$HH�� �#  H�H�hH�L$8H��$�   H��$�   H��$�   H�$H�T$`H�T$H�l$hH�l$H��$�   H�\$�    H�T$(�\$ �� ��   H��$�   L��$�   H��L9���   H��H�H�l$`H�+H�l$h�=     ugH�kH��H�T$(H�D$HH�L$8H��H��H�l$0H9��,���H��$�   H9�w(L��$�   L��$   H��$  H��$  H���   ��    L�CL�$H�l$�    H�T$(��    냉 �����H�\$@H�� tH�K H�L$pH�{(H�|$x�7�����������L�B(L�$H�D$�    H�T$@�����������    ��'���H�$H�l$L�    L�D$�    � �����    ����������������
      �  ,type.*go/ast.ValueSpec   �   "".copyConstType   � (runtime.writeBarrier   �  $"".hasExportedName   �
  ."".(*reader).filterSpec   � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �   type.go/ast.Spec   �  (runtime.panicdottype   �  0runtime.morestack_noctxt   ��  ,"".autotmp_0524   type.go/ast.Spec "".autotmp_0523  "type.*go/ast.Spec "".autotmp_0522  type.int "".autotmp_0521  type.int "".autotmp_0519 � type.go/ast.Spec "".autotmp_0518 �"type.*go/ast.Spec "".autotmp_0517 �type.int "".autotmp_0516 �type.int "".autotmp_0515  $type.[]go/ast.Spec "".autotmp_0513  type.bool "".autotmp_0512  $type.[]go/ast.Spec "".autotmp_0510  type.go/ast.Expr "".autotmp_0509 /$type.[]go/ast.Spec "".s � type.go/ast.Spec "".j �type.int "".spec �,type.*go/ast.ValueSpec "".spec � type.go/ast.Spec "".prevType � type.go/ast.Expr "".~r2 P$type.[]go/ast.Spec "".tok @&type.go/token.Token "".list $type.[]go/ast.Spec "".r  type.*"".reader "������ � ��9x#�?sE=<		 ( ���JF Tgclocals·d8668e205667c6ef4f74e27331326ebc Tgclocals·e127204208a449a4bc3afdf4417ef9c1   :$GOROOT/src/go/doc/exports.go�."".(*reader).filterDecl  �  �dH�%    H;a��  H��pH��$�   H��$�   H�L$HH�$H�D$PH�D$�    H�|$HH�t$P�T$���~�ueH��1�H9�tH�[H�-    H9��V  H��H��   < t9H�YH�� t+H�kH�M H�$H�MH�L$�    �\$��$�   H��pÉ�с���f[��   H��1�H9�tH�[H�-    H9���   H��H��   �� ��   H�\$xH�$H�� ��   H�X H�|$H�H�H�KH�OH�KH�OH�D$@H�hH�l$ �    H�T$(H�L$0H�D$8H�\$@H�� tRH�L$`H�K(H�D$hH�C0H�T$X�=     uH�S H�\$@H�k(H�� ��$�   H��p�L�C L�$H�T$�    �҉몉 �W���Ƅ$�    H��p�1�1��%���1�1������    �$�������
      v  $runtime.ifacethash   �  *type.*go/ast.FuncDecl   �  "go/ast.IsExported   �  (type.*go/ast.GenDecl   �  6"".(*reader).filterSpecList   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   @�  "".autotmp_0529 O type.go/ast.Decl "".autotmp_0528  type.bool "".autotmp_0526 /$type.[]go/ast.Spec "".d _(type.*go/ast.GenDecl "".~r1 0type.bool "".decl  type.go/ast.Decl "".r  type.*"".reader :�������+��� � 6�j9=�  :f�� Tgclocals·f7aa1743939cae014f83a8a2d262049c Tgclocals·d3b071704863cbd459bbd46f550e3b94   :$GOROOT/src/go/doc/exports.go�0"".(*reader).fileExports  �  �dH�%    H�D$�H;A��  H��   1�H�t$ H��$�   H�� �n  H�SH�C H�k(H��$�   1�H��$�   H�D$(H�T$xH��H�l$(H9���   H�D$8H�� �  H�H�hH�L$0H�T$PH�l$XH��$�   H�$H�T$@H�T$H�l$HH�l$�    H�t$ �\$�� ��   H��$�   H�� ��   H�KH�C H�k(H�l$pH��H�L$`H��H�D$hH9���   H��H�H�l$@H�+H�l$H�=     uOH�kH��H�t$ H�D$8H�L$0H��H��H�l$(H9�����H��$�   L�C(L9�wH�s H�Đ   ��    L�CL�$H�l$�    H�t$ ��    ��C���딉 �����������    �I������������
      �  ."".(*reader).filterDecl   � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt    �  "".autotmp_0538  type.go/ast.Decl "".autotmp_0537 �"type.*go/ast.Decl "".autotmp_0536 �type.int "".autotmp_0535 �type.int "".autotmp_0532 /$type.[]go/ast.Decl "".d � type.go/ast.Decl "".j �type.int "".src "type.*go/ast.File "".r  type.*"".reader  ����>� � @�p8]  ��1 Tgclocals·7e902992778eda5f91d29a3f0c115aee Tgclocals·9d98f0d067a7d5c31416a70b02745cb5   :$GOROOT/src/go/doc/exports.go�"".matchFields  �  �dH�%    H;a�B  H��xH��$�   1�H9��  H��H�� �  H�pH�@H�kH�l$p1�H�D$hH�D$(H�t$`H�l$(H9���   H�t$@H�H�|$0H�� ��   H�SH�CH�kH�l$X1�H�D$PH�D$H�T$HH��H�l$H9�}pH�D$8H�(H�L$ H�� tH�]H�H�$H�KH�L$H��$�   H���H�|$0H�t$@�\$�� tƄ$�   H��x�H�D$8H�L$ H��H��H�l$H9�|�H��H��H�l$(H9��5���Ƅ$�    H��xÉE �y�����0���� ������    �����
      �       �  0runtime.morestack_noctxt   0�  "".autotmp_0549 &type.**go/ast.Ident "".autotmp_0548 �type.int "".autotmp_0547 �type.int "".autotmp_0545 o&type.**go/ast.Field "".autotmp_0544 �type.int "".autotmp_0543 �type.int "".autotmp_0541 _(type.[]*go/ast.Ident "".autotmp_0540 /(type.[]*go/ast.Field "".~r2  type.bool "".f type."".Filter "".fields  ,type.*go/ast.FieldList ,����<��� � 6JF;  �� Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·7b90e273048a3c2d112e626ee7e85da5   8$GOROOT/src/go/doc/filter.go�"".matchDecl  �  �dH�%    H�D$�H;A��  H��   H��$�   H�� �~  H�K H�C(H�k0H��$�   1�H��$�   H�D$(H��$�   H��H�l$(H9��U  H�D$HH�� �,  H�H�hH�T$0H�L$PH�l$XH�L$pH�$H�l$xH�l$�    H�|$pH�t$x�T$��Z�v3�  H��1�H9�tH�[H�-    H9���  H��H��   < ��   H�� ��   H�QH�AH�iH��$�   1�H��$�   H�D$H��$�   H��H�l$H9�}mH�D$@H�(H�L$ H�� ��   H�]H�H�$H�KH�L$H��$�   H����\$�� tƄ$�   H�İ   �H�D$@H�L$ H��H��H�l$H9�|�H�D$HH�T$0H��H��H�l$(H9������Ƅ$�    H�İ   ÉE �s��������������u�H��1�H9�tH�[H�-    H9���  H��H��   < t�H�L$8H�YH�� �g  H�kH�M H�$H�MH�L$H��$�   H����\$�� tƄ$�   H�İ   �H�\$8H�� �  H�KH�kH�L$`H�$H�l$hH�l$�    L��$�   H�|$`H�t$h�T$��Bj	�u^H��1�H9�tH�[H�-    H9���   H��H��   �� t1H�hH�,$L�D$�    �\$�� tƄ$�   H�İ   �������=�O������H��1�H9�tH�[H�-    H9�uDH��H��   �� �[���H�hH�,$L�D$�    �\$�� tƄ$�   H�İ   ��*���1�1���1�1��Q��������������1�1��r���1�1��D���� �������{����    �@���
      �  $runtime.ifacethash   �  ,type.*go/ast.ValueSpec   �       �  *type.*go/ast.TypeSpec   �	       �
  $runtime.ifacethash   �  .type.*go/ast.StructType   �  "".matchFields   �  4type.*go/ast.InterfaceType   �  "".matchFields   �  0runtime.morestack_noctxt   0�  ("".autotmp_0570  type.uint32 "".autotmp_0569  type.bool "".autotmp_0568 � type.go/ast.Expr "".autotmp_0566 �&type.**go/ast.Ident "".autotmp_0565 �type.int "".autotmp_0564 �type.int "".autotmp_0561   type.go/ast.Spec "".autotmp_0560  type.go/ast.Spec "".autotmp_0559 �"type.*go/ast.Spec "".autotmp_0558 �type.int "".autotmp_0557 �type.int "".autotmp_0556  type.bool "".autotmp_0554  type.bool "".autotmp_0552 _(type.[]*go/ast.Ident "".autotmp_0551 /$type.[]go/ast.Spec "".v �*type.*go/ast.TypeSpec "".d � type.go/ast.Spec "".~r2  type.bool "".f type."".Filter "".d  (type.*go/ast.GenDecl T����I��������i��B�
 � n2ilO50'4?z9%
 " ���F]� Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 Tgclocals·8fe27e4ff3724ff01c209913c795c44d   8$GOROOT/src/go/doc/filter.go�"".filterValues  �  �dH�%    H;a�7  H��X1�H��$�   H��$�   H��$�   1�H�t$H�T$`H�D$hH�\$pH�\$P1�H�D$HH�D$ H�T$@H��H�l$ H9���   H�D$8H�(H�L$(H�l$0H�m(H�,$H�\$xH�\$�    H�t$�\$�� ��   H�\$`L�D$hL9���   H��H�l$0�=     u]H�+H��H�t$H�D$8H�L$(H��H��H�l$ H9��u���H�l$pH9�w"L�D$`L��$�   H��$�   H��$�   H��X��    H�$H�l$�    H�t$��    ��    ����������������
      �  "".matchDecl   � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   p�  "".autotmp_0577 ?type.**"".Value "".autotmp_0576 otype.int "".autotmp_0575 _type.int "".autotmp_0574   type.[]*"".Value "".autotmp_0571 / type.[]*"".Value 
"".vd Otype.*"".Value "".w type.int "".~r2 @ type.[]*"".Value "".f 0type."".Filter "".a   type.[]*"".Value  ����%� � 6j1C/(3  �� Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0   8$GOROOT/src/go/doc/filter.go�"".filterFuncs  �  �dH�%    H;a�P  H��X1�H��$�   H��$�   H��$�   1�H�t$H�T$`H�D$hH�\$pH�\$P1�H�D$HH�D$ H�T$@H��H�l$ H9���   H�D$8H�(H�L$(H�l$0H�� ��   H�]H�H�$H�KH�L$H�T$xH���H�t$�\$�� ��   H�\$`L�D$hL9���   H��H�l$0�=     u]H�+H��H�t$H�D$8H�L$(H��H��H�l$ H9��d���H�l$pH9�w"L�D$`L��$�   H��$�   H��$�   H��X��    H�$H�l$�    H�t$��    됉E �'����    �������
      �       � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   p�  "".autotmp_0585 ?type.**"".Func "".autotmp_0584 otype.int "".autotmp_0583 _type.int "".autotmp_0582  type.[]*"".Func "".autotmp_0579 /type.[]*"".Func 
"".fd Otype.*"".Func "".w type.int "".~r2 @type.[]*"".Func "".f 0type."".Filter "".a  type.[]*"".Func  ����-� � <�1C@(3  �� Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0   8$GOROOT/src/go/doc/filter.go�"".filterTypes  �  �dH�%    H�D$�H;A�M  H��   1�H��$�   H��$�   H��$�   H�D$8    H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$HH��$�   H��H�l$HH9���   H�D$`H�(H�L$PH�D$@    H�l$XH�m H�,$H��$�   H�\$�    H�D$X�\$�� ��   H��   H�� ~;H��$�   H�l$8L��$�   L9���   H��=     upH�H�\$8H��H�\$8H�D$`H�L$PH��H��H�l$HH9��Q���H�\$8H��$�   H9�w(L��$�   L��$�   H��$�   H��$�   H�İ   ��    H�$H�D$�    ��    H�� ��  H�X(H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H�\$XH�� �o  H��$�   H�K0H��$�   H�C8H��$�   �=     �+  H�S(H�t$XH�� �  H�^@H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H�\$XH�� ��  H��$�   H�KHH��$�   H�CPH��$�   �=     �y  H�S@H�t$XH�� �_  H�^XH�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H�\$XH�� �  H�L$pH�K`H�D$xH�ChH�T$h�=     ��   H�SXH�t$XH�� ��   H�^pH�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�D$XH�t$ H�T$(H�L$0H�� tiH�T$pH�PxH�L$xH���   H�t$h�=     u-H�ppL�D$@H�X0H�pHH�P`H�HxH�H�H�L�H������L�@pL�$H�t$�    H�D$X뾉 듉�C���L�CXL�$H�T$�    ���������������L�C@L�$H�T$�    �t�����<���������L�C(L�$H�T$�    ����������� �6����    �����&
      �  "".matchDecl   � (runtime.writeBarrier   �  $runtime.panicslice   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  "".filterValues   � (runtime.writeBarrier   �	  "".filterValues   �
 (runtime.writeBarrier   �  "".filterFuncs   � (runtime.writeBarrier   �  "".filterFuncs   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   p�   "".autotmp_0602 �type.**"".Type "".autotmp_0601 �type.int "".autotmp_0600 �type.int "".autotmp_0599  type.[]*"".Type "".autotmp_0598  type.int "".autotmp_0592  type.[]*"".Func "".autotmp_0591 �type.[]*"".Func "".autotmp_0590   type.[]*"".Value "".autotmp_0589 _ type.[]*"".Value "".autotmp_0587 /type.[]*"".Type "".n �type.int 
"".td �type.*"".Type "".w �type.int "".~r2 @type.[]*"".Type "".f 0type."".Filter "".a  type.[]*"".Type "������ � ��9	U	2."A���$   ��;� Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc Tgclocals·e61e23fa553179df29e88d2b566c0cc1   8$GOROOT/src/go/doc/filter.go�("".(*Package).Filter  �  �dH�%    H;a�
  H��   H��$�   H�� ��  H���   H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H��$�   H�� ��  H�L$pH���   H�D$xH���   H�T$h�=     �L  H���   H��$�   H�� �,  H���   H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H��$�   H�� ��  H�L$pH���   H�D$xH���   H�T$h�=     ��  H���   H��$�   H�� �n  H���   H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H��$�   H�� �  H�L$XH���   H�D$`H���   H�T$P�=     ��   H���   H��$�   H�� ��   H���   H�H�$H�KH�L$H�KH�L$H��$�   H�\$�    H�T$ H�L$(H�D$0H��$�   H�� t]H�L$@H���   H�D$HH���   H�T$8�=     u H���   H��$�   1�H�+H�kH�Ā   �L���   L�$H�T$�    �Љ량�I���L���   L�$H�T$�    ���������������L���   L�$H�T$�    �_�����'���������L���   L�$H�T$�    ������i���������    ��������������
      �  "".filterValues   � (runtime.writeBarrier   �  "".filterValues   � (runtime.writeBarrier   �  "".filterTypes   � (runtime.writeBarrier   �  "".filterFuncs   �	 (runtime.writeBarrier   �
  .runtime.writebarrierptr   �
  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".autotmp_0607 �type.[]*"".Func "".autotmp_0606 _type.[]*"".Type "".autotmp_0605   type.[]*"".Value "".autotmp_0604 / type.[]*"".Value "".f type."".Filter "".p   type.*"".Package "������ � \�����  Y� Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6 Tgclocals·6d07ab0a37c299682f1d85b92cb6cfd1   8$GOROOT/src/go/doc/filter.go�"".recvString  �  �dH�%    H;a�v  H��X1�H�\$pH�\$xH�L$`H�D$hH�L$8H�$H�D$@H�D$�    H�|$8H�t$@�T$��Ns;/uMH��1�H9�tH�[H�-    H9��  H��H��   < t!H�� tH�iH�l$pH�iH�l$xH��XÉ���Ø4���   H��1�H9�tH�[H�-    H9���   H��H��   �� t|H�� trH�XH�H�$H�KH�L$�    H�L$H�D$H�$    H�    H�\$H�D$   H�L$HH�L$H�D$PH�D$ �    H�\$(H�\$pH�\$0H�\$xH��XÉ �H�    H�\$pH�D$x   H��X�1�1��\���1�1�������    �m����������������
      �  $runtime.ifacethash   �  $type.*go/ast.Ident   �  *type.*go/ast.StarExpr   �  "".recvString   �  go.string."*"   �  *runtime.concatstring2   �  &go.string."BADRECV"   �  0runtime.morestack_noctxt   @�  "".autotmp_0609 ? type.go/ast.Expr "".autotmp_0608 type.string "".~r1  type.string "".recv   type.go/ast.Expr :���������� � ":#d!9|  @�� Tgclocals·aefd16b155593f6f07980a05b297ad1f Tgclocals·bade3c5f6d433f8d8fecc50019bf4c85   8$GOROOT/src/go/doc/reader.go� "".methodSet.set  �  �dH�%    H�D$�H;A�D  H��   H��$�   H�kH�� �  H�MH�EH�L$XH�D$`H�    H�$H��$�   H�\$H�L$xH�L$H��$�   H�D$�    H��$�   H�\$ H�1�H9�tH�XH�� tH�Ġ   �1�H�\$HH�\$PH�Y1�H9���   1�H��H�iH�� �z  H�}H��$�   H�MH�]H��$�   H��$�   H���G  H�� �6  H�/H�� �!  H�u H�U(H�t$8H�4$H�T$@H�T$�    H��$�   H�\$H�\$HH�\$H�\$PH�\$XH�\$hH�\$`H�\$pH�)H�,$�    H�\$H�\$xH�\$H��$�   H�    H�$�    H�D$H��H�� ��  W�H����    H�D$0H��$�   H�hH�l$x�=     �>  H�(H�l$`H�hH�l$X�=     �  H�hH�� ��   H��$�   �=     ��   H�h H�l$PH�h0H�l$H�=     ��   H�h(H�l$PH�h@H�l$H�=     uOH�h8H�D$(H�    H�$H��$�   H�\$H�\$hH�\$H�\$(H�\$�    H��$�   1�H�+H�Ġ   �L�@8L�$H�l$�    H�D$0�L�@(L�$H�l$�    H�D$0�e���L�@ L�$H�l$�    H�D$0�*���� �
���L�@L�$H�l$�    H�D$0�����H�$H�l$�    H�D$0����� �t����E ������    ������E �~����E ������    ��������������,
      �  "type."".methodSet   �  4runtime.mapaccess1_faststr   �  "".recvString   �  6go/ast.(*CommentGroup).Text   �  type."".Func   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �	 (runtime.writeBarrier   �	  "type."".methodSet   �
  $runtime.mapassign1   �
  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt    �  "".autotmp_0618  type.*"".Func "".autotmp_0617 �type.*"".Func "".autotmp_0616  type.string "".autotmp_0615 otype.string "".autotmp_0613 �type.*"".Func "".autotmp_0612 Otype.string "".list /(type.[]*go/ast.Field "".typ � type.go/ast.Expr "".recv �type.string "".name �type.string "".f *type.*go/ast.FuncDecl "".mset  "type."".methodSet 0��������� � dV_<4#�6z * v�'�'W0 Tgclocals·cebf12d22eea72c192e5960fe2f61bf0 Tgclocals·c479f047767b723c63a86ea32fdba623   8$GOROOT/src/go/doc/reader.go� "".methodSet.add  �  �dH�%    H;a��  H��8H�    H�$H�\$@H�\$H�t$HH�� ��  H�^H�|$H�H�H�KH�O�    H�L$HH�\$ H�1�H9��  H�YHH�hHH9���   1�H9���   H�YHH�hHH9���   H�    H�$�    H�D$H��H�� ��   W�H����    H�\$HH�� ��   H�kH�D$0L�@L�D$H�l$H�-    H�,$�    H�L$HH�D$0H�� tRH�iHH�hHH�D$(H�    H�$H�\$@H�\$H�L$H�|$ tH�D$H�\$(H�\$�    H��8É%    �݉ 몉�l���� �J���H�L$(H�    H�$H�\$@H�\$H�L$H�|$ tH�D$H�\$(H�\$�    H��8É%    �݉�v����    �1����
      4  "type."".methodSet   �  4runtime.mapaccess1_faststr   �  type."".Func   �  "runtime.newobject   ��  runtime.duffzero   �  type.string   �  (runtime.typedmemmove   �  "type."".methodSet   �  $runtime.mapassign1   �  "type."".methodSet   �  $runtime.mapassign1   �  0runtime.morestack_noctxt    p  "".autotmp_0622  type.*"".Func "".autotmp_0621  type.*"".Func "".autotmp_0620 type.*"".Func "".autotmp_0619 type.*"".Func "".m type.*"".Func "".mset  "type."".methodSet  p�op[opo � L�M.@<	<	  R�T� Tgclocals·7e902992778eda5f91d29a3f0c115aee Tgclocals·008e235a1392cc90d1ed9ad2f7e76d87   8$GOROOT/src/go/doc/reader.go�"".baseTypeName  �  �dH�%    H;a��  H��81��D$` 1�H�\$PH�\$XH�L$@H�D$HH�L$(H�$H�D$0H�D$�    H�|$(H�t$0�L$��Ns;/uRH��1�H9�tH�[H�-    H9��T  H��H��   < t&H�� tH�jH�l$PH�jH�l$X�D$` H��8É�����+�e��   H��1�H9�tH�[H�-    H9���   H��H��   �� tbH��H�(E1�L9�tH�mL�    L9�u@H�kH��   �� t+H�hH�� tH�]H�\$PH�]H�\$X�D$`H��8ÉE ��H��8�1��ǁ�Ø4�u�H��1�H9�tH�[H�-    H9�uTH��H��   �� t�H�� t;H�XH�H�$H�KH�L$�    H�L$H�D$�\$ H�L$PH�D$X�\$`H��8É ��1�1��1�1�����1�1������    �������������
      �  $runtime.ifacethash   �  $type.*go/ast.Ident   �  2type.*go/ast.SelectorExpr   �  $type.*go/ast.Ident   �  *type.*go/ast.StarExpr   �  "".baseTypeName   �  0runtime.morestack_noctxt   Pp  
"".autotmp_0625  type.go/ast.Expr "".autotmp_0624  type.bool "".imported @type.bool "".name  type.string "".x   type.go/ast.Expr 2p�op�op	opuopo � 4�*d&9.+
1E  G�V Tgclocals·ac82343006770597a842747caad5b201 Tgclocals·21a8f585a14d020f181242c5256583dc   8$GOROOT/src/go/doc/reader.go�,"".(*reader).isVisible  �  �dH�%    H;avDH��H�l$ H�] H��H�� u&H�\$(H�$H�\$0H�\$�    �\$�\$8H����D$8���    �������
      t  "go/ast.IsExported   �  0runtime.morestack_noctxt   @0  "".~r1 0type.bool "".name type.string "".r  type.*"".reader 08/0/ ` �@ 
 9' Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�."".(*reader).lookupType  �  �dH�%    H;a�  H��   H��$�   H�� tCH��uQH��$�   H�,$H�D$H�-    H�l$H�D$   �    H��$�   �\$ �� tHǄ$�       H�Ā   �H��$�   H�    H�$H��$�   H�k`H�l$H�L$pH�L$H�D$xH�D$�    H�D$ �\$(H�(�� tH��$�   H�Ā   �H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$XH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$PH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$HH�    H�$�    H�|$H��H�� ��  W�H����    H�D$8H��$�   H�hH��$�   �=     �7  H�hH�� �"  H�l$X�=     ��   H�h0H�� ��   H�l$P�=     ��   H�hPH�� ��   H�l$H�=     urH�hXH��$�   H�\$`H��$�   H�\$hH�D$0H�D$@H�    H�$H��$�   H�k`H�l$H�\$`H�\$H�\$@H�\$�    H�\$0H��$�   H�Ā   �L�@XL�$H�l$�    H�D$8�v���� �]���L�@PL�$H�l$�    H�D$8�7���� ����L�@0L�$H�l$�    H�D$8������ �����L�@L�$H�l$�    H�D$8������t����    ����������������2
      �  go.string."_"   �   runtime.eqstring   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".namedType   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �	  :type.map[string]*"".namedType   �
  $runtime.mapassign1   �
  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   @�  "".autotmp_0636 �$type.*"".namedType "".autotmp_0634 $type.*"".namedType "".autotmp_0633 ?type.string "".autotmp_0632 o"type."".methodSet "".autotmp_0631 _"type."".methodSet "".autotmp_0630 O&type."".embeddedSet "".autotmp_0629 type.string "".typ �$type.*"".namedType "".~r1 0$type.*"".namedType "".name type.string "".r  type.*"".reader :�d��^������� � >�"IO
55�Yp . T�5�
'###+ Tgclocals·573eebd23f15bbede97c85018d63627a Tgclocals·39612780d40568a5b01933408425e52c   8$GOROOT/src/go/doc/reader.go�B"".(*reader).recordAnonymousField  �  �dH�%    H�D$�H;A��  H��   1�1�H��$�   H��$�   H��$�   H�$H��$�   H�\$�    H�L$H��$�   H�T$H��$�   �\$ H��H��$�   1�H9���  < �|  H��$�   H�\$@H�L$pH��H�T$xH�� tEH����   H�$H�D$H�-    H�l$H�D$   �    H�L$pH�D$x�\$ �� ��   1�1�H9�twH��   @�h(H��$�   1�H9�tH�[H�-    H9�uUH��$�   H��   H�D$P�L$7H�    H�$H��$�   H�k0H�l$H�\$PH�\$H�\$7H�\$�    H�Ġ   �1��H�    H�$H�\$@H�k`H�l$H��$�   H�L$H��$�   H�D$�    H�D$ �\$(H�(�� tH���$���H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$hH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$`H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$XH�    H�$�    H�|$H��H�� �q  W�H����    H�D$HH�l$xH�hH�l$p�=     �)  H�hH�� �  H�l$h�=     ��   H�h0H�� ��   H�l$`�=     ��   H�hPH�� ��   H�l$X�=     ugH�hXH�\$pH��$�   H�\$xH��$�   H�D$8H�D$PH�    H�$H�\$@H�k`H�l$H��$�   H�\$H�\$PH�\$�    H�D$8�t���L�@XL�$H�l$�    H�D$H넉 �k���L�@PL�$H�l$�    H�D$H�E���� �(���L�@0L�$H�l$�    H�D$H����� �����L�@L�$H�l$�    H�D$H���������H�Ġ   ��    ���������:
      �  "".baseTypeName   �  go.string."_"   �   runtime.eqstring   �  *type.*go/ast.StarExpr   �  &type."".embeddedSet   �  $runtime.mapassign1   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �	  runtime.makemap   �	  "type."".namedType   �	  "runtime.newobject   �
�  runtime.duffzero   �
 (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   `�   "".autotmp_0646 �$type.*"".namedType "".autotmp_0644 �type.bool "".autotmp_0643  $type.*"".namedType "".autotmp_0642 �$type.*"".namedType "".autotmp_0641 ?type.string "".autotmp_0640 �"type."".methodSet "".autotmp_0639 "type."".methodSet "".autotmp_0638 o&type."".embeddedSet "".autotmp_0637 type.string "".typ �$type.*"".namedType "".name _type.string "".r �type.*"".reader "".fname @type.string "".fieldType   type.go/ast.Expr "".parent $type.*"".namedType "".r  type.*"".reader "������ � :�3@n.>� < L��Dz5�
 ##, Tgclocals·24bdc3afac682cc4abeb732876105abc Tgclocals·e4edfcfe053f06aa2f3f9df5ba415e02   8$GOROOT/src/go/doc/reader.go�("".(*reader).readDoc  �  �dH�%    H;a�  H��xH��$�   H�$�    H��$�   H�t$H�T$H�XH�� u4H�T$PH�PH�t$H�=     u	H�pH��x�L�@L�$H�t$�    ��H�HH�hH�$    H�L$hH�L$H�l$pH�l$H�    H�\$H�D$    H�t$HH�t$(H�T$PH�T$0�    H�L$8H�D$@H��$�   H�� t4H�D$`H�CH�L$X�=     u	H�KH��x�L�CL�$H�L$�    �����    �����������������
      H  6go/ast.(*CommentGroup).Text   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  go.string."\n"   �  *runtime.concatstring3   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".autotmp_0647 type.string "".text _type.string "".comment 2type.*go/ast.CommentGroup "".r  type.*"".reader ,�L������ � :�#
�  #� Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6 Tgclocals·709a14768fab2805a378215c02f0d27f   8$GOROOT/src/go/doc/reader.go�*"".(*reader).remember  �  �dH�%    H;a��   H��PH�\$XH�SxH���   H���   H��H��H9�w1H���   H��H�l$`�=     uH�+H��P�H�$H�l$�    ��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�D$0H�L$8H�\$XH�� tQH��H�D$@H��H���   H���   H�T$H�=     u	H�Sx�h���L�CxL�$H�T$�    H�T$HH�D$@�G������    ��������������
      � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  8type.[]*go/ast.InterfaceType   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".typ 4type.*go/ast.InterfaceType "".r  type.*"".reader  �B���� � "�>�  c�+ Tgclocals·2f2d69f12d345ece4be5273d9b84f0bb Tgclocals·0c8aa8e80191a30eac23f1a218103f16   8$GOROOT/src/go/doc/reader.go�"".specNames  �  �dH�%    H�D$�H;A��  H���   1�H��$  H��$  H��$  H��$�   H�    H�$H�D$    H�D$�    L�\$L��$�   L�T$ L��$�   L�L$(L��$�   H��$�   H��$�   H��$   H��$�   H�D$X    H��$�   H�D$PH��$�   H�L$hH�\$XH�l$PH9��Q  H�\$hH�� �$  H�+H�CH��$�   H��$�   H�D$xH�l$pE1�L9�tH�mL�    L9���  H��H�� ��  H�pH�@H�kH��$�   1�H��$�   H�D$@H��$�   H�l$@H9���   H�t$`H�H�|$HH�� �`  H�kH��$�   H�kH��$�   L��L��L��H��L9���   I��H��$�   H��H��Hk�H�H��$�   H�kH��$�   �=     ufH�+H��H��H�l$@H9��o���H�\$hH��H�\$hH�\$XH��H�\$XH�\$XH�l$PH9������L��$  L��$  L��$  H���   �H�$H�l$�    L��$�   L��$�   L��$�   H�|$HH�t$`�h���H�-    H�,$H�L$H�D$L�L$H�\$ �    H�|$HH�t$`L�\$(L�T$0L�L$8L��I��L��$�   L��$�   L��L��$�   ����������� �B���H�,$L�D$L�    L�L$�    �������    �����
      �  type.[]string   �  "runtime.makeslice   �  ,type.*go/ast.ValueSpec   � (runtime.writeBarrier   �	  .runtime.writebarrierptr   �
  type.[]string   �
  "runtime.growslice   �   type.go/ast.Spec   �  (runtime.panicdottype   �  0runtime.morestack_noctxt   `�  "".autotmp_0663 �type.string "".autotmp_0661 �&type.**go/ast.Ident "".autotmp_0660 �type.int "".autotmp_0659 �type.int "".autotmp_0658 � type.go/ast.Spec "".autotmp_0657 �"type.*go/ast.Spec "".autotmp_0656 �type.int "".autotmp_0655  type.int "".autotmp_0654 _(type.[]*go/ast.Ident "".autotmp_0653 /$type.[]go/ast.Spec "".autotmp_0652 �type.int "".s � type.go/ast.Spec "".names �type.[]string "".~r1 0type.[]string "".specs  $type.[]go/ast.Spec "������
 � >�9M�to. 0j#
  Z�Kg Tgclocals·adb3347b296419e60da36d67f8b7ce43 Tgclocals·a4ac9012e8051c074b7cac5858bd5519   8$GOROOT/src/go/doc/reader.go�,"".(*reader).readValue  �%  �%dH�%    H��$ ���H;A�=	  H��  1�H��$  I��H��$  H�D$H    1�H��$�   I��H��$�   H�D$@    H��$�  H�� ��  L�K H�C(H�k0H��$x  E1�H��$p  H�D$XL��$h  H�l$XI9�}|L��$�   I�� ��  I�I�AL�T$`H��$   H��$(  H��$�   H��$�   1�H9�tH�[H�-    H9��A  H��H��   < ��  I��I��H�l$XI9�|�H�\$@H�� uH�Ā  �H��$�  H�� �m  H��HH�D$hH��$  H�� �M  H��$�  H�$L�\$H�T$�    �\$�� �$  H��$�  H�[(H�l$H�H*�f(��    �Y��H,�H9���  H��$�  H�\$xH��$  H��$�   H��$  H��$�   H�� tKH����  H�$H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� ��  1�1�H9�tH�� ��  H��8H�D$hH��$�  H�+H�,$�    H�\$H��$@  H�\$H��$H  H��$�  H�� �G  H�^ H�H�$H�KH�L$H�KH�L$�    H�\$H��$P  H�\$ H��$X  H�\$(H��$`  H�\$hH�kH�l$`H�    H�$�    H�D$H��$�   H��$H  H�hH��$@  �=     ��  H�(H��$X  H�hH��$`  H�h H��$P  �=     �H  H�hH�� �3  H��$�  �=     ��   H�h(H�l$`H�h0H��$�   H�\$hH�H�kH�KH��H��H9�wAH�kH��H��$�   �=     uH�+H��$�  1�H�+H�Ā  �H�$H�l$�    ��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�l$0H�L$8H�\$hH�� tLH��H�l$PH��H�kH�KH��$�   �=     uH��Y���H�$H�T$�    H��$�   H�D$P�9�����L�@(L�$H�l$�    H��$�   ������ �����L�@L�$H�l$�    H��$�   ����H�$H�l$�    H��$�   �Q��������� �b���H�    H�$H�\$xH�k`H�l$H��$@  H�L$H��$H  H�D$�    H�D$ �\$(H�(�� tH�������H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H�    H�$�    H�|$H��H�� ��  W�H����    H��$�   H��$�   H�hH��$�   �=     �J  H�hH�� �5  H��$�   �=     �  H�h0H�� ��   H��$�   �=     ��   H�hPH�� ��   H��$�   �=     usH�hXH��$�   H��$0  H��$�   H��$8  H�D$pH��$�   H�    H�$H�\$xH�k`H�l$H��$0  H�\$H��$�   H�\$�    H�D$p�(���L�@XL�$H�l$�    H��$�   �r���� �V���L�@PL�$H�l$�    H��$�   �-���� ����L�@0L�$H�l$�    H��$�   ������ �����L�@L�$H�l$�    H��$�   ������[�������� ����1�H��$�   H��H��$�   H�i H�� �9  H�Y H�H�$H�KH�L$�    L��$  L�T$`L��$�   H��$�   H��$  H��$�   H�t$H��$   H�l$H��$  �\$ �� uH��H��$�   H��H�� tyH�� tPH��$�   H9���   L�$H�T$H�|$H�D$�    L�T$`L��$�   H��$�   H��$�   �\$ �� tSI��H��$  H��H��$  H�\$HH��H�\$HI��H��$�   H��$�   H��H��$�   H�\$@H��H�\$@����1�H��$  I������H��$�  H�]H��@�)���L��L��$�   H������1�1������A��g���������    ������������������\
      �  ,type.*go/ast.ValueSpec   �  ,"".(*reader).isVisible   �  *$f64.3fe8000000000000   �  go.string."_"   �   runtime.eqstring   �	  6go/ast.(*CommentGroup).Text   �
  "".specNames   �  type."".Value   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �   type.[]*"".Value   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".namedType   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  "".baseTypeName   �"   runtime.eqstring   �%  0runtime.morestack_noctxt    �  @"".autotmp_0689 �type.*"".Value "".autotmp_0688  type.*"".Value "".autotmp_0687 �$type.*"".namedType "".autotmp_0685 � type.go/ast.Spec "".autotmp_0684 �"type.*go/ast.Spec "".autotmp_0683 �type.int "".autotmp_0682 �type.int "".autotmp_0681  type.int "".autotmp_0680 _type.[]string "".autotmp_0679  type.string "".autotmp_0678 �$type.*"".namedType "".autotmp_0677 �type.string "".autotmp_0676 �"type."".methodSet "".autotmp_0675 �"type."".methodSet "".autotmp_0674 �&type."".embeddedSet "".autotmp_0673 type.string "".autotmp_0672  type.int "".autotmp_0670  type.int "".autotmp_0667 /$type.[]go/ast.Spec "".typ �$type.*"".namedType "".name �type.string "".r �type.*"".reader "".values �"type.*[]*"".Value "".n �type.string "".name �type.string "".spec � type.go/ast.Spec "".n �type.int "".prev �type.string "".domFreq �type.int "".domName �type.string "".decl (type.*go/ast.GenDecl "".r  type.*"".reader 0"��������
� � ��"
		~-Fo�
.[�?�`�EjV=0-
#	 f ��NNE�&"T(AS}8�
&&&\�� Tgclocals·696dc48efaf7c9921882eba1b5b5885e Tgclocals·f76a807c7b8b6a371ade38b5b9694ecd   8$GOROOT/src/go/doc/reader.go�"".fields  �  �dH�%    H;a�  H��01��D$` 1�H�\$HH�\$PH�\$XH�D$    H�L$8H�D$@H�L$ H�$H�D$(H�D$�    L�D$ H�|$(H�t$�T$��Bj	�ufL��1�I9�tH�[H�-    H9���   H��H��   < t:H�q�D$`1�H9�t!H�� t H�nH�l$HH�nH�l$PH�nH�l$XH��0É�܁�=�O�u�L��1�I9�tH�[H�-    H9�uH��H��   �� t�H�p�1�1���1�1��|����    ����������

      �  $runtime.ifacethash   �  .type.*go/ast.StructType   �  4type.*go/ast.InterfaceType   �  0runtime.morestack_noctxt   ``  
"".autotmp_0693  type.go/ast.Expr "".fields /,type.*go/ast.FieldList "".isStruct Ptype.bool "".list  (type.[]*go/ast.Field "".typ   type.go/ast.Expr `�_`J_ � <�/	i!1
  U� Tgclocals·f86cabb45f3736e32e1652a4ce443e9b Tgclocals·368ff6680f3872f8e014b9f8c1a308ff   8$GOROOT/src/go/doc/reader.go�*"".(*reader).readType  �  �dH�%    H�D$�H;A�D  H���   H��$�   H�\$PH��$   H�kH�� �  H�MH��$�   H�EH��$�   H�� tKH���J  H�$H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� �	  1�1�H9�uH���   �H�D$HH�� ��  H��$�   �=     ��  H�h H��$   H�H��$   1�H�+1�H9�uH��$�   H�H��$�   1�H�+H�$�    H�L$H�D$H�\$HH�� �R  H��$�   H�CH��$�   �=     �  H�1�H��$�   H��$�   H��$�   H��$   H�� ��   H�^H�H�$H�KH�L$�    H�L$H�D$H�T$ H�\$H�l$(@�k)H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$0H��$�   H��H�l$0H9�}dH�T$XH�H�t$8H�hH�� uUH��$�   H�$H�\$HH�\$H�X H�|$H�H�H�KH�O�    H�t$8H�T$XH��H��H�l$0H9�|�H���   �������H�$H�L$�    ����������L�@ L�$H�l$�    �7���� ����H�    H�$H�\$PH�k`H�l$H��$�   H�L$H��$�   H�D$�    H�D$ �\$(H�(�� tH������H�    H�$H�D$    H�D$    H�D$    �    H�\$ H��$�   H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$xH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$pH�    H�$�    H�|$H��H�� ��  W�H����    H�D$`H��$�   H�hH��$�   �=     �5  H�hH�� �   H��$�   �=     ��   H�h0H�� ��   H�l$x�=     ��   H�hPH�� ��   H�l$p�=     umH�hXH��$�   H��$�   H��$�   H��$�   H�D$@H�D$hH�    H�$H�\$PH�k`H�l$H��$�   H�\$H�\$hH�\$�    H�D$@�����L�@XL�$H�l$�    H�D$`�{���� �b���L�@PL�$H�l$�    H�D$`�<���� ����L�@0L�$H�l$�    H�D$`������ �����L�@L�$H�l$�    H�D$`������v����E ������    ��������������@
      �  go.string."_"   �   runtime.eqstring   � (runtime.writeBarrier   �  6go/ast.(*CommentGroup).Text   � (runtime.writeBarrier   �  "".fields   �	  B"".(*reader).recordAnonymousField   �
  .runtime.writebarrierptr   �
  .runtime.writebarrierptr   �
  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".namedType   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   0�  ("".autotmp_0709 �&type.**go/ast.Field "".autotmp_0708 �type.int "".autotmp_0707 �type.int "".autotmp_0706 �$type.*"".namedType "".autotmp_0703 /(type.[]*go/ast.Field "".autotmp_0702  type.string "".autotmp_0701 �$type.*"".namedType "".autotmp_0700 �type.string "".autotmp_0699 �"type."".methodSet "".autotmp_0698 �"type."".methodSet "".autotmp_0697 �&type."".embeddedSet "".autotmp_0696 type.string "".typ �$type.*"".namedType "".name �type.string "".r �type.*"".reader "".list _(type.[]*go/ast.Field "".typ �$type.*"".namedType "".spec  *type.*go/ast.TypeSpec "".decl (type.*go/ast.GenDecl "".r  type.*"".reader 0��������� �
 ���
(F
HQ
<
	
	M�� B ���:b}5�
###2 Tgclocals·e76d9788ffeb8eb69a0d7b2c884b94ed Tgclocals·7301d8fdff8300440e17cffa48be7961   8$GOROOT/src/go/doc/reader.go�*"".(*reader).readFunc  �"  �"dH�%    H�D$�H;A�Z  H���   H��$   1�H�h H�X1�H9���  H�hH�� ��  H�MH�EH�]H��$�   H��$�   H�� H��$�   ��  H�H�� �n  H�k H�M H�$H�MH�L$�    H�L$H�T$�\$ �� tH���   �H��$�   H�\$@H�L$xH��$�   H��$�   H��H��$�   H�� tCH��uhH�$H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� t+1�1�H9�tH�hXH�,$H��$   H�\$�    H���   �H�    H�$H�\$@H�k`H�l$H��$�   H�L$H��$�   H�D$�    H�D$ �\$(H�(�� tH���H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$pH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$hH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$`H�    H�$�    H�|$H��H�� ��  W�H����    H�D$PH��$�   H�hH��$�   �=     �2  H�hH�� �  H�l$p�=     ��   H�h0H�� ��   H�l$h�=     ��   H�hPH�� ��   H�l$`�=     umH�hXH��$�   H��$�   H��$�   H��$�   H�D$0H�D$XH�    H�$H�\$@H�k`H�l$H��$�   H�\$H�\$XH�\$�    H�D$0�����L�@XL�$H�l$�    H�D$P�{���� �b���L�@PL�$H�l$�    H�D$P�<���� ����L�@0L�$H�l$�    H�D$P������ �����L�@L�$H�l$�    H�D$P������y���������    �E �A���H�XH�kH�,$�    H�\$H���D  H��$   H�kH�]H�� �#  H�KH�CH�kH��$�   H��$�   H�� H��$�   ��  H�H�hH����  H�X H�H�$H�KH�L$�    H�T$H��$�   H�L$H��$�   �\$ �� ��  H��$�   H�$H�T$H�L$�    �\$�� �i  H��$�   H�\$HH��$�   H��$�   H��$�   H��$�   H�� tGH����   H�$H�D$H�-    H�l$H�D$   �    H��$�   H��$�   �\$ �� tU1�1�H9�t"H�hPH�,$H��$   H�\$�    H���   �H��$�   H�khH�,$H��$   H�\$�    H���   �H�    H�$H�\$HH�k`H�l$H��$�   H�L$H��$�   H�D$�    H�D$ �\$(H�(�� tH���[���H�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$pH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$hH�    H�$H�D$    H�D$    H�D$    �    H�\$ H�\$`H�    H�$�    H�|$H��H�� ��  W�H����    H�D$PH��$�   H�hH��$�   �=     �2  H�hH�� �  H�l$p�=     ��   H�h0H�� ��   H�l$h�=     ��   H�hPH�� ��   H�l$`�=     umH�hXH��$�   H��$�   H��$�   H��$�   H�D$8H�D$XH�    H�$H�\$HH�k`H�l$H��$�   H�\$H�\$XH�\$�    H�D$8����L�@XL�$H�l$�    H�D$P�{���� �b���L�@PL�$H�l$�    H�D$P�<���� ����L�@0L�$H�l$�    H�D$P������ �����L�@L�$H�l$�    H�D$P������y����7����2����    �����������    ��������r
      �  "".baseTypeName   �  go.string."_"   �   runtime.eqstring   �   "".methodSet.set   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �	  "type."".namedType   �	  "runtime.newobject   �	�  runtime.duffzero   �
 (runtime.writeBarrier   �
 (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  :go/ast.(*FieldList).NumFields   �  "".baseTypeName   �  ,"".(*reader).isVisible   �  go.string."_"   �   runtime.eqstring   �   "".methodSet.set   �   "".methodSet.set   �  :type.map[string]*"".namedType   �  4runtime.mapaccess2_faststr   �  &type."".embeddedSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".methodSet   �  runtime.makemap   �  "type."".namedType   �  "runtime.newobject   ��  runtime.duffzero   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �   .runtime.writebarrierptr   �!  .runtime.writebarrierptr   �!  $runtime.panicindex   �!  0runtime.morestack_noctxt    �  2"".autotmp_0729  $type.*"".namedType "".autotmp_0728  &type.**"".namedType "".autotmp_0727 �$type.*"".namedType "".autotmp_0725  $type.*"".namedType "".autotmp_0724  type.string "".autotmp_0723  "type."".methodSet "".autotmp_0722  "type."".methodSet "".autotmp_0721  &type."".embeddedSet "".autotmp_0720  type.string "".autotmp_0716 �$type.*"".namedType "".autotmp_0715 otype.string "".autotmp_0714 �"type."".methodSet "".autotmp_0713 �"type."".methodSet "".autotmp_0712 �&type."".embeddedSet "".autotmp_0711 Otype.string "".typ �$type.*"".namedType "".name �type.string "".r �type.*"".reader "".typ �$type.*"".namedType "".name �type.string "".r �type.*"".reader "".n �type.string "".recvTypeName �type.string "".fun *type.*go/ast.FuncDecl "".r  type.*"".reader J����������)���� � n�'r�$ Kj�"�
 S v �x=@w5�
###	�n=jz5�
### ! Tgclocals·715f4247ff054ce54b6559cd80f93589 Tgclocals·e7cc1a3a5ad7e5bd5d4932eddee30345   8$GOROOT/src/go/doc/reader.go�*"".(*reader).readNote  �  �dH�%    H��$h���H;A��  H��  1�H��$�   H��$�   H��$�   H��$�   H��$(  H�(H��$0  H�hH��$8  H�hH�$�    H�L$H�D$H�    H�$H�L$XH�L$H�D$`H�D$�    H�D$H�L$ H�\$(H��$�   H�� �@  H��H��$�   H��H��$�   ��  H��H�H�l$`H9���  L�D$XH)�H�� tM�L��$�   L�$H��$�   H�l$H�D$   �    H��$�   H��$�   H�\$H�\$xH�D$ H��$�   H�� ��  H��H���W  H��H�H��H���<  H��H�+L�D$`L9��   H9��  L�D$XH)�H�� tM�L��$�   H��$�   L�D$hH�l$pH��H�    H�$H��$   H�k0H�l$L��$�   L�D$H��$�   H�L$�    H��$(  H��$�   H��$�   H��$0  H�\$ H�� �w  H�+H��$   H�kH��$  H�kH��$  H�� �C  H�/H�m H�l$HH��H��H9��!  H�,�H�E H�HH�H�H�\$@H��H����  H�� H�H��H����  H��(H�+L�D$`L9���  H9���  L�D$XH)�H�� tM� H��$�   L��$�   H�    H�$�    H�D$H�l$HH�(H�l$@H�hH�D$PH��$�   H�hH��$�   �=     �,  H�hH��$�   H�h(H�l$x�=     ��   H�h H�D$PH��$   H��$  H��$  H��H��H9���   H��H��H��$�   H��$�   H��$�   H��H�l$P�=     uFH�+H�    H�$H��$   H�k0H�l$H��$�   H�\$H��$�   H�\$�    H��  �H�$H�l$�    �H�-    H�,$H�T$H�D$H�L$H�\$ �    H�T$(H�D$0H�L$8�B���L�@ L�$H�l$�    H�D$P�����L�@L�$H�l$�    H�D$P�����    �    �    �    �    ������    �    �    �    �    �    �"�����<
      �  6go/ast.(*CommentGroup).Text   �  "".noteMarkerRx   �  Pregexp.(*Regexp).FindStringSubmatchIndex   �  "".clean   �  4type.map[string][]*"".Note   �  4runtime.mapaccess1_faststr   �  type."".Note   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  4type.map[string][]*"".Note   �  $runtime.mapassign1   �  .runtime.writebarrierptr   �  type.[]*"".Note   �  "runtime.growslice   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   @�  ,"".autotmp_0749 �type.*"".Note "".autotmp_0748  type.*"".Note "".autotmp_0746 �0type.go/ast.CommentGroup "".autotmp_0744 _type.[]*"".Note "".autotmp_0743 �type.string "".autotmp_0742  type.int "".autotmp_0741  type.int "".autotmp_0740  type.int "".autotmp_0739  type.int "".autotmp_0738 /type.[]*"".Note "".autotmp_0737  type.string "".autotmp_0736 �type.string "".autotmp_0734  type.int "".autotmp_0733 �type.string "".~r0 �"type.go/token.Pos "".~r0 �"type.go/token.Pos "".marker �type.string "".body �type.string "".m �type.[]int "".text �type.string "".list ,type.[]*go/ast.Comment "".r  type.*"".reader ""������ �	 r�"XE
�Q�&aU�H : k.����<&*/ Tgclocals·d40c6564e2ba8bed9102651873b34d14 Tgclocals·bddc76d8a57f9840df311eb725104ff2   8$GOROOT/src/go/doc/reader.go�,"".(*reader).readNotes  �
  �
dH�%    H�D$�H;A�  H���   H��$�   H��$�   H��$�   H��$�   H�D$H    H��$�   H�D$@H��$�   H�L$XH�\$HH�l$@H9���  H�\$XH�H������H�L$(H�� ��  H�;H�kH�l$hH�sH�|$`H�T$hH�t$pH��$�   1�H��$�   H�T$0H��$�   H��H�l$0H9���   H�T$PH�*H�D$8H�D$ H�    H�$H�� �  H�]H�|$H�H�H�KH�O�    H�|$`H�t$pH�L$(�\$�� �A  H�� |lH�l$ I��H9��#  H9��  H)�I)�I��I�� tM��H��$�   H�$L�L$xL�L$H��$�   H�l$L��$�   L�D$�    H�|$`H�t$pH�L$ H�L$(H�T$PH�D$8H��H��H�l$0H9�����H�� |\H�l$hI��H9���   H)�I)�I��I�� tM��H��$�   H�$L��$�   L�L$H��$�   H�l$L��$�   L�D$�    H�\$XH��H�\$XH�\$HH��H�\$HH�\$HH�l$@H9�����H���   ��    �    �6����E �y����������    �_������������������
      �   "".noteCommentRx   �  8regexp.(*Regexp).MatchString   �  *"".(*reader).readNote   �  *"".(*reader).readNote   �	  $runtime.panicslice   �	  $runtime.panicslice   �
  0runtime.morestack_noctxt   @�  "".autotmp_0764 �*type.**go/ast.Comment "".autotmp_0763 �type.int "".autotmp_0762 �type.int "".autotmp_0760 �4type.**go/ast.CommentGroup "".autotmp_0759 �type.int "".autotmp_0758 �type.int "".autotmp_0757  ,type.[]*go/ast.Comment "".autotmp_0756 �,type.[]*go/ast.Comment "".autotmp_0754 _,type.[]*go/ast.Comment "".autotmp_0753 /6type.[]*go/ast.CommentGroup "".j �type.int "".list �,type.[]*go/ast.Comment "".i �type.int "".comments 6type.[]*go/ast.CommentGroup "".r  type.*"".reader  ����"� � T�^QNl
	\.  ��;; Tgclocals·14c16763214c88f6ebc22b4b638329b7 Tgclocals·db3311d7e1cb6ec5029186017096a081   8$GOROOT/src/go/doc/reader.go�*"".(*reader).readFile  �!  �!dH�%    H��$���H;A�  H��p  H��$�  H�] 1�H9�t.H��$x  H�$H��$�  H�+H�l$�    H��$�  1�H�+H��$�  H�� ��  H�KH�C H�k(H��$h  1�H��$`  H�D$HH��$X  H��H�l$HH9���   H��$�   H�� �^  H�H�hH�T$PH��$�   H��$�   H��$  H�$H��$  H�l$�    H��$  H��$  �T$���~���   H��1�H9�tH�[H�-    H9���  H��H��   < ��   H��$x  H�$H�L$�    H��$�   H�T$PH��H��H�l$HH9��,���H��$x  H�$H��$�  H�� tBH�^hH�|$H�H�H�KH�OH�KH�O�    H��$�  1�H�khH�kpH�kxH��p  É뺁���f[�r���H��1�H9�tH�[H�-    H9��   H��H��   �� �A���H�hH��K�a  H��@uH��$x  H�$H�D$�    ����H��K����H��H�H H�@(H�k0H��$P  H�D$@    H��$H  H�D$8H��$@  H��$�   H�\$@H�l$8H9������H��$�   H�� ��  H�H�CH��$�   H��$   H��$�   H��H��$�   1�H9�tH�[H�-    H9��  H��H��   < �8  H�L$`H�YH�� �S  H�kH�M H�$H�MH�L$�    H�T$H��$�   H�L$H��$�   H�D$ H�\$(H��$�   H��$�   H�� ��   H��$  H��$   H�D$X   H�    H�$H��$x  H�k8H�l$H��$  H�\$H�\$XH�\$�    H�D$`H�X1�H9�tlH�hH�� ��   H�MH��$�   H�EH��$�   H��u@H�$H�D$H�-    H�l$H�D$   �    �\$ �� tH��$x  H��   @�k@H��$�   H��H��$�   H�\$@H��H�\$@�&����E �t��������1�1�������,���H��T�e  H�h(H����   H�hH�� ���� ��   H�X H�H(H�h0H��$P  H��$@  H�� H��$H  vUH�+E1�L9�tH�mL�    L9�u4H�SH��   �� �M���H��$x  H�$H�D$H�T$�    �-���1�1����    H��H�D$pH�� ��  H�P H�@(H�k0H��$P  1�H��$H  H�D$8H��$@  H�l$8H9������H��$�   H�� �R  H�H�BH�t$@H��$�   H��$   H��$�   H��$�   1�H9�tH�[H�-    H9��  H��H��   < �h  H�iH�m H�l$0H�L$hH��$�   H�    H�$�    H�D$1�H�(H�hH�hH�hH�h H�h(H�h0H�h8H�D$xH�l$pL�E �=     �m  L� H�l$0H�hH�@T   H�    H�$�    H�\$H�� �3  HǄ$0     HǄ$8     H��$(  H�    1�H9���   H��$�   H��$(  H��$�   H�H��$   �=     ��   H�KH�\$xH��$0  H�k(H��$8  H�k0H��$(  �=     uBH�k H�D$xH��$x  H�$H�D$H�\$hH�\$�    H�t$@H��$�   H��H������L�C L�$H�l$�    �L�CL�$H�L$�    �e���H�    H�$H�    H�\$H�    H�\$�    H�D$�����������H�$L�D$�    H�D$x�~���1�1������������ �U���H��U�,����T���1�1�����1�1��$���� ������F����    ������������F
      �  ("".(*reader).readDoc   �  $runtime.ifacethash   �  *type.*go/ast.FuncDecl   �  *"".(*reader).readFunc   �  ,"".(*reader).readNotes   �  (type.*go/ast.GenDecl   �	  ,"".(*reader).readValue   �  .type.*go/ast.ImportSpec   �  strconv.Unquote   �  &type.map[string]int   �  $runtime.mapassign1   �  go.string."."   �   runtime.eqstring   �  *type.*go/ast.TypeSpec   �  *"".(*reader).readType   �  $runtime.panicindex   �  *type.*go/ast.TypeSpec   �  &type.go/ast.GenDecl   �  "runtime.newobject   � (runtime.writeBarrier   �  &type.[1]go/ast.Spec   �  "runtime.newobject   �  Hgo.itab.*go/ast.TypeSpec.go/ast.Spec   � (runtime.writeBarrier   � (runtime.writeBarrier   �  *"".(*reader).readType   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  *type.*go/ast.TypeSpec   �   type.go/ast.Spec   �  Hgo.itab.*go/ast.TypeSpec.go/ast.Spec   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �   0runtime.morestack_noctxt    �  H"".autotmp_0796 �$type.[]go/ast.Spec "".autotmp_0795 �(type.*go/ast.GenDecl "".autotmp_0793   type.go/ast.Spec "".autotmp_0792  "type.*go/ast.Spec "".autotmp_0791  type.int "".autotmp_0790  type.int "".autotmp_0788 �type.string "".autotmp_0787 � type.go/ast.Spec "".autotmp_0786 �"type.*go/ast.Spec "".autotmp_0785 �type.int "".autotmp_0784 �type.int "".autotmp_0780   type.go/ast.Decl "".autotmp_0779 � type.go/ast.Decl "".autotmp_0778 �"type.*go/ast.Decl "".autotmp_0777 �type.int "".autotmp_0776 �type.int "".autotmp_0775  *type.*go/ast.TypeSpec "".autotmp_0774  *type.*go/ast.TypeSpec "".autotmp_0773  $type.[]go/ast.Spec "".autotmp_0772 �*type.*go/ast.TypeSpec "".autotmp_0771  type.int "".autotmp_0770 �type.int "".autotmp_0769 �type.string "".autotmp_0767 _$type.[]go/ast.Spec "".autotmp_0766 /$type.[]go/ast.Decl "".~r0 �"type.go/token.Pos "".s �*type.*go/ast.TypeSpec "".spec � type.go/ast.Spec "".err �type.error "".import_ �type.string "".s �.type.*go/ast.ImportSpec "".spec � type.go/ast.Spec "".d �(type.*go/ast.GenDecl "".decl � type.go/ast.Decl "".src "type.*go/ast.File "".r  type.*"".reader ""������ � ��"!l~jk"v>s=#
�8kVd	&	
"Y76
�5C�-!P	
 X Q�f`���_��e�+-f Tgclocals·a21ab7bae19632fedab25371b764faba Tgclocals·3eb79ea418853034459ea0e413208728   8$GOROOT/src/go/doc/reader.go�0"".(*reader).readPackage  �  �dH�%    H�D$�H;A�(  H��   H��$  H�] 1�H9�tH�H��H�    H�$H�D$H�D$�    H�T$H�L$ H�D$(H��$  H�� ��  H��$�   H�K H��$�   H�C(H��$�   �=     ��  H�SH�    H�$H�D$    H�D$    H�D$    �    H�D$ H��$  H�� �5  �=     �  H�C8H��$  H��$  H�+H�    H�$H�D$    H�D$    H�D$    �    H�D$ H��$  H�� ��  �=     ��  H�C`H�    H�$H�D$    H�D$    H�D$    �    H�D$ H��$  H�� �@  �=     �  H�ChH�    H�$H�D$    H�D$    H�D$    �    H�D$ H��$  H�� ��  �=     ��  H�C0H�D$0    H��$  H�k H��$�   W�H����    H�    H�$H�l$H��$�   H�\$�    H��$�   1�H9���   H��$�   H�� �0  H�H�CH��$  H�� �  H�sH�S H�k(H��$�   H��H��$�   H�l$0H��$�   H9���  H��H�H�D$pH�CH�L$h�=     ��  H�H�\$0H��H�\$0H��$�   H�$�    H��$�   1�H9��J���H��$  H�� �R  H�^H�H�$H�KH�L$H�KH�L$�    H��$  H�� �  H�KH�C H�k(H��$�   1�H��$�   H�D$8H��$�   H��H�l$8H9���   H�D$PH�� ��   H�H�@H�T$@H�L$XH�D$`H�    H�$H��$  H�k H�l$H�L$xH�L$H��$�   H�D$�    H�\$ H�H��$  H��H�� u H��$  H�$H�D$HH�D$�    H�D$HH��$  H�$H�D$�    H�D$PH�T$@H��H��H�l$8H9��4���H��   É �4��������������H�$H�L$�    �Q����    ������������L�C0L�$H�D$�    �B�����*���L�ChL�$H�D$�    ����������L�C`L�$H�D$�    �`�����H���L�C8L�$H�D$�    �����������L�CL�$H�T$�    �k�����3����    ����������D
      v  type.[]string   �  "runtime.makeslice   � (runtime.writeBarrier   �  &type.map[string]int   �  runtime.makemap   � (runtime.writeBarrier   �  :type.map[string]*"".namedType   �  runtime.makemap   � (runtime.writeBarrier   �  "type."".methodSet   �  runtime.makemap   � (runtime.writeBarrier   �  4type.map[string][]*"".Note   �  runtime.makemap   � (runtime.writeBarrier   ��  runtime.duffzero   �  8type.map[string]*go/ast.File   �	  &runtime.mapiterinit   � (runtime.writeBarrier   �  &runtime.mapiternext   �  sort.Strings   �  8type.map[string]*go/ast.File   �  4runtime.mapaccess1_faststr   �  0"".(*reader).fileExports   �  *"".(*reader).readFile   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   0�  """.autotmp_0817 �type.string "".autotmp_0816 �type.*string "".autotmp_0815 �type.int "".autotmp_0814  type.int "".autotmp_0812  type.string "".autotmp_0811  type.[]string "".autotmp_0810  type.int "".autotmp_0809 �Btype.map.iter[string]*go/ast.File "".autotmp_0803 �type.[]string "".autotmp_0802 �type.int "".f �"type.*go/ast.File "".filename �type.string "".filename �type.string "".i �type.int "".mode  type."".Mode "".pkg (type.*go/ast.Package "".r  type.*"".reader "������ �
 ���SSSS	nl$4iJ 		 . M���5J,� Tgclocals·42e7756549fd1f1e78e70fcb9f08dd2b Tgclocals·7fe2912721285589731dc5ce1f08c6a7   8$GOROOT/src/go/doc/reader.go� "".customizeRecv  �  �dH�%    H�D$�H;A�?  H��   H��$�   1�H9��  H�X 1�H9��  H�h H�]1�H9���  H�h H�]H�kH����  H�    H�$�    H�T$H��$�   H�k H�]H�� ��  H�KH�CH�kH��$�   H��$�   H�� H��$�   �r  H�)H�� �]  H�T$XH�T$H�l$H�-    H�,$�    H�\$XH�K H�k(H��$�   H�,$H�L$xH�Y(��H�\$H�\$(H�\$XH�k E1�L9�tH�mL�    L9���  H�k(�D$'H�    H�$�    H�D$1�H�(H�hH�hH�hH�l$(H�(H�D$@H��$�   H�hH��$�   �=     �h  H�hH��H�D$0H�D$@H�    1�H9��  H�T$@H�T$pH�D$h��$�    ��   �|$' ��   H�)H��H�)H�L$@H�    H�$�    H�T$H�T$8H�l$(H�*H�    1�H9��m  H�L$@H�� �W  H�D$xH�BH��$�   �=     �  H�JH�T$8H�    1�H9���  H�T$8H�\$XH�D$hH�C H�T$p�=     ��  H�S(H�    H�$�    H�D$H��$�   H�k H�]H�� �Z  H�D$PH�D$H�\$H�    H�$�    H�    H�$�    H�D$H�� �  HǄ$�      HǄ$�      H��$�   H�l$X�=     ��  H�(H�\$PH��$�   H�kH��$�   H�k�=     ��  H�CH�    H�$�    H�D$H��$�   H�k H�� �M  H�D$HH�D$H�l$H�-    H�,$�    H�\$HH�l$P�=     �   H�kH�    H�$�    H�D$H��$�   H�� ��   H�D$`H�D$H�\$H�    H�$�    H�\$`H�l$H�=     ��   H�k H�\$hH�$H�\$pH�\$�    H�T$`H�L$H�D$H��$�   H�B0H��$�   �=     u H�J(H��$�   H�jHH��$�   H�İ   �L�B(L�$H�L$�    H�T$`��L�C L�$H�l$�    �l�����+���L�CL�$H�l$�    ������E ����L�CL�$H�D$�    �i���H�$H�l$�    H��$�   � ���� ����������L�C(L�$H�T$�    �Y���H�    H�$H�    H�\$H�    H�\$�    H�D$�����L�BL�$H�L$�    H�T$8����������H�    H�$H�    H�\$H�    H�\$�    H�T$8H�D$�\���H�    H�$H�    H�\$H�    H�\$�    H�L$0H�D$����L�@L�$H�l$�    H�D$@�����D$' �����E �����    ��R���H��$�   H�İ   ��    �������������������v
      �  "type.go/ast.Field   �  "runtime.newobject   �  "type.go/ast.Field   �  (runtime.typedmemmove   �       �  *type.*go/ast.StarExpr   �  "type.go/ast.Ident   �  "runtime.newobject   � (runtime.writeBarrier   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �  (type.go/ast.StarExpr   �  "runtime.newobject   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �	 (runtime.writeBarrier   �	  Hgo.itab.*go/ast.StarExpr.go/ast.Expr   �
 (runtime.writeBarrier   �
  *type.go/ast.FieldList   �
  "runtime.newobject   �  *type.go/ast.FieldList   �  (runtime.typedmemmove   �  *type.[1]*go/ast.Field   �  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   �  (type.go/ast.FuncDecl   �  "runtime.newobject   �  (type.go/ast.FuncDecl   �  (runtime.typedmemmove   � (runtime.writeBarrier   �  type."".Func   �  "runtime.newobject   �  type."".Func   �  (runtime.typedmemmove   � (runtime.writeBarrier   �  "".recvString   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  *type.*go/ast.StarExpr   �   type.go/ast.Expr   �  Hgo.itab.*go/ast.StarExpr.go/ast.Expr   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  $type.*go/ast.Ident   �   type.go/ast.Expr   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �   runtime.typ2Itab   �  $type.*go/ast.Ident   �   type.go/ast.Expr   �  Bgo.itab.*go/ast.Ident.go/ast.Expr   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   `�  ,"".autotmp_0830  (type.[]*go/ast.Field "".autotmp_0829  type.*uint8 "".autotmp_0828  type.*uint8 "".autotmp_0827 �*type.*go/ast.StarExpr "".autotmp_0825 �$type.*go/ast.Ident "".autotmp_0824 Otype.string "".autotmp_0823  *type.*go/ast.StarExpr "".autotmp_0822  $type.*go/ast.Ident "".autotmp_0820  $type.*go/ast.Ident "".&newField �$type.*go/ast.Field  "".&newFieldList �,type.*go/ast.FieldList "".&newFuncDecl �*type.*go/ast.FuncDecl "".&newF �type.*"".Func "".typ � type.go/ast.Expr "".newIdent �$type.*go/ast.Ident  "".origRecvIsPtr �type.bool "".origPos �"type.go/token.Pos "".~r4 Ptype.*"".Func "".level @type.int  "".embeddedIsPtr 0type.bool "".recvTypeName type.string "".f  type.*"".Func "������ � ��'C
�..[+	�$N�JFH"	�7 \ uy��>�:+63w--U7!!7 Tgclocals·86c3de611c79526d490a82204ab8e699 Tgclocals·705a498ed8ccdac9185f030fb45a87b7   8$GOROOT/src/go/doc/reader.go�F"".(*reader).collectEmbeddedMethods  �  �dH�%    H��$H���H;A�~  H��8  H��$P  H�\$p�D$GH�    H�$H��$x  H�\$H�\$pH�\$H�\$GH�\$�    H��$P  H�k0H��$�   W�H����    H�    H�$H�l$H��$�   H�\$�    H��$�   1�H9��  H��$�   �+H��$�   H���$h   ��  @�l$FH�L$XH�iXH�|$xW�H����    H�    H�$H�l$H�\$xH�\$�    H�\$x1�H9���  H��$�   H�H�\$xH�� �B  H�XHH�� ��  H��$H  H�\$HH�$H��$X  H�\$H��$`  H�\$�\$F�\$H��$p  H�\$ �    H�D$(H�    H�$H�\$HH�\$H�D$PH�� ��  H�XH�|$H�H�H�KH�O�    H�L$PH�\$ H�1�H9��@  H�YHH�hHH9��/  1�H9���   H�YHH�hHH9���   H�    H�$�    H�|$H��H�� ��  W�H����    H�\$PH�� ��  H�kH�D$`H�� ��  L�@L�D$H�l$H�-    H�,$�    H�L$`H�D$PH�� �u  H�hHH�iHH�L$hH�    H�$H�\$HH�\$H�D$H�|$ �6  H�D$H�\$hH�\$�    H�\$xH�$�    H�\$x1�H9�� ���H�D$XH�    H�$H��$x  H�\$H�D$�    H�\$�+@�� ��   H��$@  H�$H��$H  H�\$H�\$XH�\$H��$X  H�\$H��$`  H�\$ �\$F�\$(H��$p  H��H�\$0H��$x  H�\$8�    H��$�   H�$�    H��$�   1�H9������H��$P  H�\$pH�    H�$H��$x  H�\$H�\$pH�\$�    H��8  �랉%    ���������� �K�����1��������H�L$hH�    H�$H�\$HH�\$H�L$H�|$ tH�D$H�\$hH�\$�    �v����%    �݉ �;���������D$F�J����    �]����������������:
      n  &type."".embeddedSet   �  $runtime.mapassign1   ��  runtime.duffzero   �  &type."".embeddedSet   �  &runtime.mapiterinit   ��  runtime.duffzero   �  "type."".methodSet   �  &runtime.mapiterinit   �   "".customizeRecv   �  "type."".methodSet   �  4runtime.mapaccess1_faststr   �  type."".Func   �  "runtime.newobject   �	�  runtime.duffzero   �
  type.string   �
  (runtime.typedmemmove   �
  "type."".methodSet   �  $runtime.mapassign1   �  &runtime.mapiternext   �  &type."".embeddedSet   �  2runtime.mapaccess1_fast64   �  F"".(*reader).collectEmbeddedMethods   �  &runtime.mapiternext   �  &type."".embeddedSet   �  "runtime.mapdelete   �  "type."".methodSet   �  $runtime.mapassign1   �  0runtime.morestack_noctxt   ��  ."".autotmp_0853  type.*"".Func "".autotmp_0852 �type.*"".Func "".autotmp_0850  $type.*"".namedType "".autotmp_0849  type.bool "".autotmp_0847  type.*"".Func "".autotmp_0846 �type.*"".Func "".autotmp_0845  type.*"".Func "".autotmp_0844  type.*"".Func "".autotmp_0843 �:type.map.iter[string]*"".Func "".autotmp_0841 �@type.map.iter[*"".namedType]bool "".autotmp_0839 �type.bool "".autotmp_0838 �$type.*"".namedType "".m �type.*"".Func "".mset �"type."".methodSet ("".thisEmbeddedIsPtr �type.bool "".embedded �$type.*"".namedType "".visited p&type."".embeddedSet "".level `type.int  "".embeddedIsPtr Ptype.bool "".recvTypeName 0type.string "".typ  $type.*"".namedType "".mset "type."".methodSet "".r  type.*"".reader ""������ �	 ^�	"Ckc�9h$"4#d 8 `Bu~E�\7
zXnB Tgclocals·11c63aa4b444ca1a56e95d01623cf60d Tgclocals·ff840c582379ce333f10594801100e10   8$GOROOT/src/go/doc/reader.go�<"".(*reader).computeMethodSets  �	  �	dH�%    H��$ ���H;A�/  H��`  W�H�|$x�    G�H��$h  H�k`H��$   W�H����    H�    H�$H�l$H��$   H�\$�    H��$   1�H9��*  H��$  H�H��$   H�� ��  H�D$P�X)�� ��   1�H�\$x��$�   ��$�   ��$�   H��$�   H��$�   H��$�   H��$�   H��$�   W�H����    G�H�    H�$H�D$    H�\$xH�\$H��$�   H�\$�    H�L$PH�D$ H��$h  H�$H�iXH�l$H�L$H�YH�|$H�H�H�KH�O�D$( H�D$0   H�D$8�    H��$   H�$�    H��$   1�H9������H��$h  �]p�� ttH��$h  H�� tnH�SxH���   H���   H�l$p1�H�D$hH�D$@H�T$`H��H�l$@H9�}1H�D$XH�(H�L$HH�,$�    H�D$XH�L$HH��H��H�l$@H9�|�H��`  É뎉�[����    ����������������
      V�  runtime.duffzero   ��  runtime.duffzero   �  :type.map[string]*"".namedType   �  &runtime.mapiterinit   ��  runtime.duffzero   �  &type."".embeddedSet   �  runtime.makemap   �  F"".(*reader).collectEmbeddedMethods   �  &runtime.mapiternext   �  &"".removeErrorField   �	  0runtime.morestack_noctxt   �  "".autotmp_0863 �6type.**go/ast.InterfaceType "".autotmp_0862 �type.int "".autotmp_0861 �type.int "".autotmp_0860 �Dtype.map.bucket[*"".namedType]bool "".autotmp_0859 �>type.map.hdr[*"".namedType]bool "".autotmp_0857 �8type.[]*go/ast.InterfaceType "".autotmp_0855 �Dtype.map.iter[string]*"".namedType "".t �$type.*"".namedType "".r  type.*"".reader  "����� � >�	3r�$P	  p�S�I Tgclocals·5d2b5a2aeff4e4cf961f497a12cc05ae Tgclocals·81bdb1fcce921ebe87bf14577379b26e   8$GOROOT/src/go/doc/reader.go�2"".(*reader).cleanupTypes  �  �dH�%    H��$����H;A��  H��  H��$�  H�k`H��$H  W�H����    H�    H�$H�l$H��$H  H�\$�    H��$H  1�H9��  H��$P  H�+H��$H  H�� �}  H��$�  H�$H�l$HH�� �Z  H�]H�|$H�H�H�KH�O�    H�L$H�\$�\$GH�Y 1�H9�uoH�    H�$H�    H�\$H�YH�|$H�H�H�KH�O�    H�L$HH�\$ �+@�� ��   �|$G t�Y(�� ��   H��$�  �]@�� u}H�Y 1�H9�t3�|$G t,H��$H  H�$�    H��$H  1�H9������H�Ĩ  �H�    H�$H��$�  H�k`H�l$H�L$H�|$ tH�D$�    랉%    ��H��$�  H�� �   H�sHL�CPH�CXH�� �  H�i8H��$�   H�y@H�iHH��$�   H��$�   L��$�   H��$�   H��L��L��$�   H��$�   H�H)�H��H�� ~[H�    H�$H��$�   H�t$L�D$H��$�   H�L$H�D$ �    L��$�   H��$�   H�t$(H�\$0H��$�   H�L$8H�    H�$L��L��H�I��H��$�   H9��   H9��  H)�I)�I��H��$�   I�� tM��H�l$L�D$L�L$H��$�   H�\$ H�|$(H��$�   H�\$0�    H��$�   H��$�   H��$�   H�H9���  H��H��$�  H�CPH�KXH��$�   �=     �_  H�kHH�\$HH�kPH��$�   W�H����    H�    H�$H�l$H��$�   H�\$�    H��$�   1�H9���   H��$�   H�H��$�   H�� ��  H�H�kH�T$`H��$�   H�l$hH��$�   H�D$XH�    H�$H��$�  H�khH�l$H��$�   H�\$H�\$XH�\$�    H��$�   H�$�    H��$�   1�H9��a���H�\$HH�kXH��$�   W�H����    H�    H�$H�l$H��$�   H�\$�    H�L$HH��$�   1�H9��   H��$�   H�H��$�   H�� ��   H�H�kH�D$PH�L$pH�l$xH��H�    H�$H��$�  H�khH�l$H��$�   H�L$H��$�   H�D$�    �\$(�� u\H�\$pH��$�   H�\$xH��$�   H�\$PH�\$XH�    H�$H��$�  H�khH�l$H��$�   H�\$H�\$XH�\$�    H��$�   H�$�    H�L$HH��$�   1�H9�� �����������������L�CHL�$H�l$�    �����    �    �������������E ������|����    �������������������D
      |�  runtime.duffzero   �  :type.map[string]*"".namedType   �  &runtime.mapiterinit   �  ,"".(*reader).isVisible   �  (type.map[string]bool   �  &"".predeclaredTypes   �  4runtime.mapaccess1_faststr   �  &runtime.mapiternext   �  :type.map[string]*"".namedType   �  "runtime.mapdelete   �	   type.[]*"".Value   �
  &runtime.growslice_n   �
  type.*"".Value   �  ,runtime.typedslicecopy   � (runtime.writeBarrier   ��  runtime.duffzero   �  "type."".methodSet   �  &runtime.mapiterinit   �  "type."".methodSet   �  $runtime.mapassign1   �  &runtime.mapiternext   ��  runtime.duffzero   �  "type."".methodSet   �  &runtime.mapiterinit   �  "type."".methodSet   �  4runtime.mapaccess2_faststr   �  "type."".methodSet   �  $runtime.mapassign1   �  &runtime.mapiternext   �  .runtime.writebarrierptr   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   �  &"".autotmp_0883  type.*"".Func "".autotmp_0880 � type.[]*"".Value "".autotmp_0879 � type.[]*"".Value "".autotmp_0878 � type.[]*"".Value "".autotmp_0876  type.*"".Func "".autotmp_0875  type.string "".autotmp_0874 �type.string "".autotmp_0873  :type.map.iter[string]*"".Func "".autotmp_0872  "type."".methodSet "".autotmp_0871 �type.*"".Func "".autotmp_0870 �type.string "".autotmp_0869 �:type.map.iter[string]*"".Func "".autotmp_0866 �Dtype.map.iter[string]*"".namedType "".m �type.*"".Func "".name �type.string "".name �type.string "".visible �type.bool "".t �$type.*"".namedType "".r  type.*"".reader ""�����	� � x�
"rEz.1$:434	!�vW$�R\) F _g������f=
C Tgclocals·a9ea41aae9e32efcc8711d8fabe405fb Tgclocals·cf6154774c0aa37b6123d9727e16ac04   8$GOROOT/src/go/doc/reader.go�"".(*data).Len      H�\$H�+H�l$���     "".~r0 type.int "".d  type.*"".data   �
  Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�"".(*data).Swap  �  �dH�%    H;av*H��H�\$ H�$H�\$(H�\$H�l$H�UH���H����    ��
      d       t  0runtime.morestack_noctxt   0   "".j  type.int "".i type.int "".d  type.*"".data  % @ �
@ 
 2 Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�"".(*data).Less  �  �dH�%    H;av3H��H�\$(H�$H�\$0H�\$H�l$ H�UH����\$�\$8H����    ��������
      d       �  0runtime.morestack_noctxt   @0  "".~r2 0type.bool "".j  type.int "".i type.int "".d  type.*"".data 0./ P �
P 
 2 Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�"".sortBy  �  �dH�%    H;a��   H��8H�    H�$�    H�D$H�l$PH�(H�D$ H�l$H�=     ��   H�hH�� ��   H�l$@�=     uhH�hH�D$ H�    1�H9�t"H�L$ H�D$(H�$H�L$0H�L$�    H��8�H�    H�$H�    H�\$H�    H�\$�    H�D$�L�@L�$H�l$�    H�D$ 냉 �j���L�@L�$H�l$�    H�D$ �D����    ����������������
      4  type."".data   F  "runtime.newobject   � (runtime.writeBarrier   � (runtime.writeBarrier   �  >go.itab.*"".data.sort.Interface   �  sort.Sort   �  type.*"".data   �  &type.sort.Interface   �  >go.itab.*"".data.sort.Interface   �   runtime.typ2Itab   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   0p  
"".autotmp_0886 /type.*"".data "".autotmp_0885  type.*"".data "".n  type.int "".swap &type.func(int, int) "".less  0type.func(int, int) bool p�opko � �
�k  "�] Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60   8$GOROOT/src/go/doc/reader.go�"".sortedKeys  �  �dH�%    H�D$�H;A��  H���   1�H��$�   H��$�   H��$�   H��$�   1�H9�tH�H��H�    H�$H�D$H�D$�    H�\$H�\$HH�\$ H�\$PH�\$(H�\$XH�D$0    H��$�   H�|$`W�H����    H�    H�$H�D$H�\$`H�\$�    H�\$`1�H9�tvH�\$`H�� ��   H�H�CH�\$HH�l$0L�D$PL9���   H��H�H�D$@H�CH�L$8�=     u{H�H�\$0H��H�\$0H�\$`H�$�    H�\$`1�H9�u�H�\$HH�$H�\$PH�\$H�\$XH�\$�    H�\$HH��$�   H�\$PH��$�   H�\$XH��$�   H���   �H�$H�L$�    �u����    ��'����    �;��������������
      �  type.[]string   �  "runtime.makeslice   ��  runtime.duffzero   �  &type.map[string]int   �  &runtime.mapiterinit   � (runtime.writeBarrier   �  &runtime.mapiternext   �  sort.Strings   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  0runtime.morestack_noctxt   @�  "".autotmp_0893  type.int "".autotmp_0892 �0type.map.iter[string]int "".key �type.string "".i �type.int "".list �type.[]string "".~r1 type.[]string "".m  &type.map[string]int  ����!� � <�
9M	Z9"/  c_�=
# Tgclocals·c87a734079562d73ffd9eee8328c7183 Tgclocals·ef5fd2c82c386cd66d746b952cc06875   8$GOROOT/src/go/doc/reader.go�"".sortingName  �  �dH�%    H;a��   H�L$1�H�i(H����   H��H�I H�C(H�k0H��H�� ��   H�)E1�L9�tH�mL�    L9�ucH�KH��   < tGH��H�� t:H�IH�CH�kH�� v!H�)H�� tH�]H�\$H�]H�\$ÉE ���    ���1�H�\$H�\$�1�1���    ���    �%��������

      �  ,type.*go/ast.ValueSpec   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0   "".~r1 type.string "".d  (type.*go/ast.GenDecl � � $�FG  �6 Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�"".sortedValues  �
  �
dH�%    H�D$�H;A�[  H��   1�H��$�   H��$�   H��$�   H��$�   H�    H�$H�D$H�D$�    H�\$H�\$`H�\$ H�\$hH�\$(H�\$p1�H��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$8H�T$xH�l$8H9�}bH�T$XH�H�t$@H�h(H�]H��$�   H9�u/H�\$`H�L$0L�D$hL9��y  H�ˀ=     �F  H�H��H��H��H�l$8H9�|�H�l$pH9��  H�L$hH�L$@H�    H�$�    H�D$H�-    H�(H�D$PH�l$hH�hH�l$pH�hH�l$`�=     ��   H�hH�    H�$�    H�D$H�-    H�(H�D$HH�l$hH�hH�l$pH�hH�l$`�=     uPH�hH�\$PH�$H�D$H�\$@H�\$�    H�\$`H��$�   H�\$hH��$�   H�\$pH��$�   H�Đ   �L�@L�$H�l$�    H�D$H�L�@L�$H�l$�    �<����    H�$H�D$�    H�t$@H�T$XH�L$0�����    �    �������&
      �   type.[]*"".Value   �  "runtime.makeslice   � (runtime.writeBarrier   �  Vtype.struct { F uintptr; list []*"".Value }   �  "runtime.newobject   �  *"".sortedValues.func1   � (runtime.writeBarrier   �  Vtype.struct { F uintptr; list []*"".Value }   �  "runtime.newobject   �  *"".sortedValues.func2   � (runtime.writeBarrier   �  "".sortBy   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �	  $runtime.panicslice   �	  .runtime.writebarrierptr   �	  $runtime.panicindex   �	  0runtime.morestack_noctxt   p�  "".autotmp_0907 �Xtype.*struct { F uintptr; list []*"".Value } "".autotmp_0906 Xtype.*struct { F uintptr; list []*"".Value } "".autotmp_0904 otype.**"".Value "".autotmp_0903 �type.int "".autotmp_0902  type.int "".autotmp_0901  type.int "".autotmp_0899 / type.[]*"".Value "".autotmp_0898 �type.int "".i �type.int "".list _ type.[]*"".Value "".~r2 @ type.[]*"".Value "".tok 0&type.go/token.Token "".m   type.[]*"".Value  ����`� � `�9@K,
LH/	 , V�LUA
 Tgclocals·4a5c83272286258cf484ac950366f973 Tgclocals·ad7181e2240ebb348baa41afdc8d0afe   8$GOROOT/src/go/doc/reader.go�"".sortedTypes  �  �dH�%    H��$@���H;A��  H��@  1�H��$X  H��$`  H��$h  H��$H  1�H9�tH�H��H�    H�$H�D$H�D$�    H�\$H�\$hH�\$ H�\$pH�\$(H�\$xH�D$8    H��$H  H��$�   W�H����    H�    H�$H�D$H��$�   H�\$�    H��$�   1�H9��U  H��$�   H�+H��$�   H�� �  H�l$HH�� ��  H�]8H�H�$H�KH�L$H�KH�L$H�D$@   �    H�\$ H��$�   H�\$(H��$�   H�\$0H��$�   H�t$HH�� ��  H�^8H�H�$H�KH�L$H�KH�L$H�D$U   �    H�\$ H��$�   H�\$(H��$�   H�\$0H��$�   H�\$HH�kPH�,$�D$�    H�\$H��$�   H�\$H��$�   H�\$ H��$�   H�\$HH�kXH�,$��$P  �\$�    H�\$H��$�   H�\$H��$�   H�\$ H��$�   H�    H�$�    H�D$H�l$HH�� ��  H�D$`H�� �|  H�D$H�l$H�-    H�,$�    H�\$HH�� �L  H�kH�\$`H�� �2  L�CL�D$H�l$H�-    H�,$�    H�\$`H�� ��  H�l$HL�E �=     ��  L�C H�\$`H��$�   H�k0H��$�   H�k8H��$�   �=     ��  H�k(H�\$`H��$�   H�kHH��$�   H�kPH��$�   �=     �7  H�k@H�\$`H��$�   H�k`H��$�   H�khH��$�   �=     ��  H�kXH�\$`H��$�   H�kxH��$�   H���   H��$�   �=     ��  H�kpH�\$hH�l$8L�D$pL9��w  H��H�l$`�=     �N  H�+H�\$8H��H�\$8H��$�   H�$�    H��$�   1�H9������H�\$pH�\$@H�    H�$�    H�D$H�-    H�(H�D$XH�l$pH�hH�l$xH�hH�l$h�=     ��   H�hH�    H�$�    H�D$H�-    H�(H�D$PH�l$pH�hH�l$xH�hH�l$h�=     uPH�hH�\$XH�$H�D$H�\$@H�\$�    H�\$hH��$X  H�\$pH��$`  H�\$xH��$h  H��@  �L�@L�$H�l$�    H�D$P�L�@L�$H�l$�    �<���H�$H�l$�    �����    L�CpL�$H�l$�    �S���L�CXL�$H�l$�    ����L�C@L�$H�l$�    ����L�C(L�$H�l$�    �i���H�k H�,$L�D$�    ���������������������� �}����E �f�����f����E ������������    ������������������T
      �  type.[]*"".Type   �  "runtime.makeslice   ��  runtime.duffzero   �  :type.map[string]*"".namedType   �  &runtime.mapiterinit   �  "".sortedValues   �  "".sortedValues   �  "".sortedFuncs   �  "".sortedFuncs   �	  type."".Type   �	  "runtime.newobject   �
  type.string   �
  (runtime.typedmemmove   �  type.string   �  (runtime.typedmemmove   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   � (runtime.writeBarrier   �  &runtime.mapiternext   �  Ttype.struct { F uintptr; list []*"".Type }   �  "runtime.newobject   �  ("".sortedTypes.func1   � (runtime.writeBarrier   �  Ttype.struct { F uintptr; list []*"".Type }   �  "runtime.newobject   �  ("".sortedTypes.func2   � (runtime.writeBarrier   �  "".sortBy   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt   P�  """.autotmp_0920 �Vtype.*struct { F uintptr; list []*"".Type } "".autotmp_0919 �Vtype.*struct { F uintptr; list []*"".Type } "".autotmp_0918 �type.*"".Type "".autotmp_0916  type.int "".autotmp_0915  type.int "".autotmp_0914 �type.[]*"".Func "".autotmp_0913 �type.[]*"".Func "".autotmp_0912 � type.[]*"".Value "".autotmp_0911 � type.[]*"".Value "".autotmp_0910 �Dtype.map.iter[string]*"".namedType "".autotmp_0908 �type.int "".t �$type.*"".namedType "".i �type.int "".list �type.[]*"".Type "".~r2  type.[]*"".Type "".allMethods type.bool "".m  :type.map[string]*"".namedType ""��	���� � ��<M	n
aa>Z8@�
1$ 
LH/	
	c	
 \ feja>E7=�-LUA
[ Tgclocals·330a8f52616cf9d268418fab976acddc Tgclocals·748e3f8a785e34acbbe52dd60e6e6e96   8$GOROOT/src/go/doc/reader.go�"".removeStar  �  �dH�%    H;av\H�L$H�D$1�H�� ~8H�� v=���*u*H��H��rH��H��H�� tH��H�l$H�\$ ��    H�L$H�D$ ��    �    ���������������
      �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   @   "".~r1  type.string "".s  type.string � � �* 
 R. Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   8$GOROOT/src/go/doc/reader.go�"".sortedFuncs  �  �dH�%    H�D$�H;A�e  H���   1�H��$  H��$  H��$  H��$�   1�H9�tH�H��H�    H�$H�D$H�D$�    H�\$H�\$xH�\$ H��$�   H�\$(H��$�   H�D$0    H��$�   H��$�   W�H����    H�    H�$H�D$H��$�   H�\$�    H��$�   1�H9�tLH��$�   H�H��$�   H�� �w  H�X 1�H9��l  H��$�   H�$�    H��$�   1�H9�u�H�\$0H��$�   H9��/  H��$�   H�\$8H�    H�$�    H�D$H�-    H�(H�D$PH��$�   H�hH��$�   H�hH�l$x�=     ��   H�hH�    H�$�    H�D$H�-    H�(H�D$HH��$�   H�hH��$�   H�hH�l$x�=     uVH�hH�\$PH�$H�D$H�\$8H�\$�    H�\$xH��$  H��$�   H��$  H��$�   H��$  H���   �L�@L�$H�l$�    H�D$H�L�@L�$H�l$�    �0����    ��$    tPH�\$xH�l$0L��$�   L9�s2H��=     uH�H�\$0H��H�\$0�Q���H�$H�D$�    ���    H�XHH�� t�H�D$@H�H8H�@@1�H�� ~mH�� vv���*u_H��H�D$pH��rJH��H��H�L$hH�� tH��H��H��H�T$XH�$H�D$`H�D$�    H�D$@�\$�� �0��������    H�L$hH��H�D$p��    ������    �y������������4
      �  type.[]*"".Func   �  "runtime.makeslice   ��  runtime.duffzero   �  "type."".methodSet   �  &runtime.mapiterinit   �  &runtime.mapiternext   �  Ttype.struct { F uintptr; list []*"".Func }   �  "runtime.newobject   �  ("".sortedFuncs.func1   � (runtime.writeBarrier   �  Ttype.struct { F uintptr; list []*"".Func }   �  "runtime.newobject   �  ("".sortedFuncs.func2   � (runtime.writeBarrier   �  "".sortBy   �	  .runtime.writebarrierptr   �	  .runtime.writebarrierptr   �	  $runtime.panicslice   �
 (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  "go/ast.IsExported   �  $runtime.panicslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   P�  "".autotmp_0933 �Vtype.*struct { F uintptr; list []*"".Func } "".autotmp_0932 �Vtype.*struct { F uintptr; list []*"".Func } "".autotmp_0930  type.int "".autotmp_0929  type.int "".autotmp_0926  type.int "".autotmp_0925 �:type.map.iter[string]*"".Func "".autotmp_0923 �type.int "".~r1 �type.string "".s �type.string "".m �type.*"".Func "".i �type.int "".list �type.[]*"".Func "".~r2  type.[]*"".Func "".allMethods type.bool "".m  "type."".methodSet "������ � ~�9S	j RN5
'�	 8 ck�R[G
	So7 Tgclocals·fb63e74b6f2618e7c5d9866e2c2934f2 Tgclocals·98894f398543f5a4f57ec3edfd994f6a   8$GOROOT/src/go/doc/reader.go�"".noteBodies  �  �dH�%    H�D$�H;A��  H��   1�H��$�   H��$�   H��$�   1�H�\$hH�\$pH�\$xH��$�   H��$�   H��$�   H��$�   1�H��$�   H�D$@H��$�   H�l$@H9���   H�t$PH�H�|$HH�� �  H�k H�l$XH�k(H�l$`H�L$hH�\$pH�T$xH��H��H9���   H�\$pH��H��Hk�H�H�l$`H�kH�l$X�=     uGH�+H��H��H�l$@H9��x���H�\$hH��$�   H�\$pH��$�   H�\$xH��$�   H�Ę   �H�$H�l$�    H�|$HH�t$P�H�-    H�,$H�L$H�D$H�T$H�\$ �    H�|$HH�t$PH�L$(H�\$0H�T$8H��H��H�\$pH�T$xH�L$h�$����������    �8�����������
      � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]string   �  "runtime.growslice   �  0runtime.morestack_noctxt   `�  "".autotmp_0939 type.string "".autotmp_0937 �type.**"".Note "".autotmp_0936 �type.int "".autotmp_0935 �type.int "".autotmp_0934 /type.[]*"".Note "".list _type.[]string "".~r1 0type.[]string "".notes  type.[]*"".Note  ����x� � ,�9Rf/^  �0Q Tgclocals·adb3347b296419e60da36d67f8b7ce43 Tgclocals·3fda2e0c42698195f82d5b8e047ca0ad   8$GOROOT/src/go/doc/reader.go�&"".firstSentenceLen  �  �dH�%    H;a�8  H��`�D$,    �D$0    �D$4    H�\$hH�\$PH�\$pH�\$X1�H�L$HH�\$PH�$H�\$XH�\$H�L$�    �l$4H�L$�D$ H�L$@H�� ��   H�\$HH�\$8��
��   ����   ��	��   �D$(�� u>��.u9�\$0�$�    �\$�� tW�\$,�$�    �l$4H�L$@�D$(�\$�� u4��0  t���  t�\$0�\$,�l$0�D$4�1���H�\$8H�\$xH��`�H�\$8H�\$xH��`ø    �l���H�\$pH�\$xH��`��    ���������������

      �  &runtime.stringiter2   �  unicode.IsUpper   �  unicode.IsUpper   �  0runtime.morestack_noctxt   0�  "".autotmp_0948 ?type.int "".autotmp_0947 /type.int "".autotmp_0946  type.int "".autotmp_0943 type.string "".q otype.int32 "".i Otype.int "".p Wtype.int32 
"".pp _type.int32 "".ppp gtype.int32 "".~r1  type.int "".s  type.string ,������� � :"^G  b� Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·d8fdd2a55187867c76648dc792366181   <$GOROOT/src/go/doc/synopsis.go�"".clean  �  �dH�%    H;a��  H��hL�\$x1�H��$�   H��$�   E1�L��M��H��    1�L9�}XH�\$pH�|$HL9��C  H�;�+H��$�   H��H��H�� �  ��
�  H��    �L$G�� uu< uqH��L9�|�H�� ~< uH��H��L9�wMH��H�$    L�T$PL�T$H�t$XH�t$L�L$`L�L$�    H�\$ H��$�   H�\$(H��$�   H��h��    L�T$PL��H�t$XH��L�L$`H��H��L9�wH��H��H���^���H�-    H�,$H�T$H�D$L�L$H�\$ �    L�\$xH�|$H�L$GL�T$(H�t$0L�L$8H��H��L��륀��������	�����������    �    �T�������
      �  2runtime.slicebytetostring   �  $runtime.panicslice   �  type.[]uint8   �  "runtime.growslice   �  $runtime.panicindex   �  0runtime.morestack_noctxt   P�  "".autotmp_0952  type.int "".autotmp_0950  type.int "".q Atype.uint8 "".i ?type.int "".b /type.[]uint8 "".~r2 0type.string "".flags  type.int "".s  type.string "������ � ^T.		
J)M  �� Tgclocals·89fe65749ce0afc971c0982226501ff0 Tgclocals·790e5cc5051fc0affc980ade09e929ec   <$GOROOT/src/go/doc/synopsis.go�"".Synopsis  �	  �	dH�%    H�D$�H;A�  H��   1�H��$�   H��$�   H��$�   H�$H��$�   H�\$�    H�\$H��$�   H9���  H��$�   H�l$pH�,$H�\$xH�\$H�D$    �    H�\$H��$�   H�\$ H��$�   H�    H�    H�    H��$�   1�H��$�   H�D$(H��$�   H��H�l$(H9���   H��H�D$8H�� �  H� H�kH�L$0H�D$pH�D$`H�l$xH�l$hH��$�   H�$H��$�   H�\$�    L�D$H�t$L�D$@H�|$`H�|$PH�D$hH�t$HH�D$XH9���   H9���   H9���   L�D$pL�$H�D$xH�D$H�|$H�D$�    �\$ H��< t1�H��$�   H��$�   H�Ę   �H�D$8H�L$0H��H��H�l$(H9�����H��$�   H��$�   H��$�   H��$�   H�Ę   �1���    1�댉 ������    �    ���������������
      �  &"".firstSentenceLen   �  "".clean   �  $"".IllegalPrefixes   � $"".IllegalPrefixes   �  $"".IllegalPrefixes   �  strings.ToLower   �   runtime.eqstring   �  $runtime.panicslice   �  $runtime.panicslice   �  0runtime.morestack_noctxt   @�  "".autotmp_0967  type.string "".autotmp_0966 �type.*string "".autotmp_0965 �type.int "".autotmp_0964  type.int "".autotmp_0963  type.string "".autotmp_0959  type.string "".autotmp_0958 /type.[]string "".autotmp_0957 Otype.string "".autotmp_0956 �type.int "strings.prefix·3 �type.string strings.s·2 �type.string "".prefix otype.string "".~r1  type.string "".s  type.string ,����F��� � 2�1ww�
(  J�ev- Tgclocals·55cc6ee7528f0b48e5a6d9bfba36524a Tgclocals·575fdb695a683406ac81277ae7ac66b5   <$GOROOT/src/go/doc/synopsis.go�"".blocks.func1  �  �dH�%    H;a�l  H��   H�ZH�\$PH�BH�\$PH�+H�� ��   1�H�\$`H�\$hH�\$pH�\$xH�D$`    H�t$PH�\$hH�H�H�NH�KH�NH�KH��H�D$XH�H�hH�HH��H��H9�wkH�kH��H��Hk� H�H�l$`H�+H�l$pH�kH�l$xH�kH�l$h�=     uH�kH�\$P1�H�+H�kH�kH�Ā   �L�CL�$H�l$�    ��H�    H�$H�T$H�D$H�L$H�l$ �    H�T$(H�D$0H�L$8H�\$XH��H�D$@H��H�kH�KH�T$H�=     uH��8���H�$H�T$�    H�T$HH�D$@�����    �w����������
      � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  type.[]"".block   �  "runtime.growslice   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  "runtime.morestack    �  "".autotmp_0969 ?type."".block "".&out O type.*[]"".block "".&para _type.*[]string "������ � *�'�~  �&K% Tgclocals·f6bd6b3389b872033d462029172c8612 Tgclocals·9edbfbd6af913bb4812a079f727a5e32   :$GOROOT/src/go/doc/comment.go�("".playExample.func1  �  �dH�%    H;a�  H��@H�|$HH�t$PH�ZH�\$8L�JL�BH�Z H�\$0H��1�H9�tH�[H�-    H9���  H��H��   < tWH�    H�$H�|$H��H�	H�H�NH�O�    H�\$H�H�$H�KH�L$H�\$8H�+H�l$�    �D$X H��@�H��1�H9�tH�[H�-    H9��3  H��H��   < tbH�    H�$H�� tMH�YH�|$H�H�H�KH�O�    H�\$H�H�$H�KH�L$H�\$8H�+H�l$�    �D$X H��@É�H��1�H9�tH�[H�-    H9���   H��H��   �� tBH�X1�H9�uJ�D$/H�    H�$L�L$H�D$H�|$ tH�D$H�\$/H�\$�    �D$XH��@É%    ��H�    H�$L�D$H�hH�l$�    H�\$�+@�� t
H�\$0���1�1��e���1�1������1�1��B����    ����������
      �  2type.*go/ast.SelectorExpr   �   type.go/ast.Node   �  runtime.convI2I   �  go/ast.Inspect   �  2type.*go/ast.KeyValueExpr   �   type.go/ast.Node   �  runtime.convI2I   �  go/ast.Inspect   �  $type.*go/ast.Ident   �  (type.map[string]bool   �  $runtime.mapassign1   �  8type.map[*go/ast.Object]bool   �  2runtime.mapaccess1_fast64   �  "runtime.morestack   0�  
"".autotmp_0976 !type.bool "".&usesTopDecl type.*bool "".&inspectFunc 8type.*func(go/ast.Node) bool "".~r1  type.bool "".n   type.go/ast.Node 2�����|�\ � T�;,M

,T
-7

		,			  �'c'�I Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 Tgclocals·008e235a1392cc90d1ed9ad2f7e76d87   :$GOROOT/src/go/doc/example.go�*"".sortedValues.func1  �  �dH�%    H�D$�H;A��  H���   H�ZH��H�H�CH�kH��$�   H9���  H��H�H�C(1�H�h(H���e  H��H�H H�@(H�k0H��$�   H��H��$�   H�� H��$�   �*  H�)E1�L9�tH�mL�    L9��  H�KH��   < ��  H��H�� ��  H�IH�CH�kH��$�   H��$�   H�� H��$�   ��  H�)H�� ��  H�uH�UH�|$(H�H�GH�oH��$�   H��$�   H��$�   H��$�   H9��?  H��H�H�C(1�H�h(H���"  H��H�H H�@(H�k0H��$�   H��H��$�   H�� H��$�   ��  H�)E1�L9�tH�mL�    L9���  H�KH��   < ��  H��H�� ��  H�IH�CH�kH��$�   H��$�   H�� H��$�   �Y  H�)H�� �D  H�MH�EH�t$0H�T$8H��H�L$@H��H�D$HH��$�   H�t$`H��$�   H��H�T$pH�T$PH�D$xH9���   H�l$`H�,$H�L$hH�L$H�l$PH�l$H�D$XH�D$�    H�T$(H�L$hH�D$X�\$ �� thH�
H�BL�BL��$�   I9�sIJ�,�H�m H�]0H�
H�BL�JL��$�   I9�sN��M� I�h0H9���$�   H���   ��    �    H�l$`H�,$H�L$hH�L$H�l$PH�l$H�D$XH�D$�    H�\$ H�� ��$�   H���   ÉE �����    ��k���1�H������1�1��C����    ���    �E �q����    ��(���1�H���a���1�1�� ����    ���    �    �+��������������
      �  ,type.*go/ast.ValueSpec   �  ,type.*go/ast.ValueSpec   �
   runtime.eqstring   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.cmpstring   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack   0�  "".autotmp_0983 �type.string "".autotmp_0982 �type.string "".autotmp_0981  ,type.*go/ast.ValueSpec "".autotmp_0980  type.int "".&list �"type.*[]*"".Value "".~r1 �type.string "".~r1 �type.string 
"".nj �type.string 
"".ni �type.string "".~r2  type.bool "".j type.int "".i  type.int ,����R��r� � �&�hEr  �x� Tgclocals·f56b2291fa344104975cb6587be42b9b Tgclocals·ce81e155410342c1a623d0fa5be5f2a2   8$GOROOT/src/go/doc/reader.go�*"".sortedValues.func2  �  �dH�%    H;a�  H��HH�t$PH�ZH��H�+H�l$0H�kH�l$8H�kH�l$@H�H�KH�kH9���   H��H�+H�l$H�H�HH�hH9���   H��H��H�H�@L�EL�D$(H�L$L�D$XH�D$ I9�siJ�,�L�E �=     uHL�H�\$0H�l$XL�D$8L9�s*H��H�l$�=     uH�+H��H�H�$H�l$�    ���    H�$L�D$�    ��    �    �    �    �����������������
      � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack    �  "".autotmp_0993 otype.*"".Value "".autotmp_0992 / type.[]*"".Value "".j type.int "".i  type.int  ����<� � 
��  �+ Tgclocals·c55cf99de9cdd8c8202a466952fa1a45 Tgclocals·f304628972275ea37e1ee36ac34113c0   8$GOROOT/src/go/doc/reader.go�("".sortedTypes.func1  �  �dH�%    H;a��   H��@H�ZH�H�KH�sH�l$HH9���   H�4�H�.H�� ��   L�EI�H�$I�HH�L$H�H�CH�sH�t$8H�L$(H�l$PH�D$0H9�sAH�4�H�.H�� t/L�EH�|$I�H�I�HH�O�    H�\$ H�� �D$XH��@ÉE ���    �E �x����    �    �"�����

      �  "runtime.cmpstring   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack   0�  "".~r2  type.bool "".j type.int "".i  type.int ��� � 
��  �? Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·790e5cc5051fc0affc980ade09e929ec   8$GOROOT/src/go/doc/reader.go�("".sortedTypes.func2  �  �dH�%    H;a�  H��HH�t$PH�ZH��H�+H�l$0H�kH�l$8H�kH�l$@H�H�KH�kH9���   H��H�+H�l$H�H�HH�hH9���   H��H��H�H�@L�EL�D$(H�L$L�D$XH�D$ I9�siJ�,�L�E �=     uHL�H�\$0H�l$XL�D$8L9�s*H��H�l$�=     uH�+H��H�H�$H�l$�    ���    H�$L�D$�    ��    �    �    �    �����������������
      � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack    �  "".autotmp_1000 otype.*"".Type "".autotmp_0999 /type.[]*"".Type "".j type.int "".i  type.int  ����<� � 
��  �+ Tgclocals·c55cf99de9cdd8c8202a466952fa1a45 Tgclocals·f304628972275ea37e1ee36ac34113c0   8$GOROOT/src/go/doc/reader.go�("".sortedFuncs.func1  �  �dH�%    H;a��   H��@H�ZH�H�KH�sH�l$HH9���   H�4�H�.H�� ��   L�EI�H�$I�HH�L$H�H�CH�sH�t$8H�L$(H�l$PH�D$0H9�sAH�4�H�.H�� t/L�EH�|$I�H�I�HH�O�    H�\$ H�� �D$XH��@ÉE ���    �E �x����    �    �"�����

      �  "runtime.cmpstring   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack   0�  "".~r2  type.bool "".j type.int "".i  type.int ��� � 
��  �? Tgclocals·790e5cc5051fc0affc980ade09e929ec Tgclocals·790e5cc5051fc0affc980ade09e929ec   8$GOROOT/src/go/doc/reader.go�("".sortedFuncs.func2  �  �dH�%    H;a�  H��HH�t$PH�ZH��H�+H�l$0H�kH�l$8H�kH�l$@H�H�KH�kH9���   H��H�+H�l$H�H�HH�hH9���   H��H��H�H�@L�EL�D$(H�L$L�D$XH�D$ I9�siJ�,�L�E �=     uHL�H�\$0H�l$XL�D$8L9�s*H��H�l$�=     uH�+H��H�H�$H�l$�    ���    H�$L�D$�    ��    �    �    �    �����������������
      � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  "runtime.morestack    �  "".autotmp_1007 otype.*"".Func "".autotmp_1006 /type.[]*"".Func "".j type.int "".i  type.int  ����<� � 
��  �+ Tgclocals·c55cf99de9cdd8c8202a466952fa1a45 Tgclocals·f304628972275ea37e1ee36ac34113c0   8$GOROOT/src/go/doc/reader.go�"".init  �  �dH�%    H;a��  H��@�    �� t�    ��uH��@��    �    �    �    �    �    �    �    �    �    �    H�    H�$H�D$�   �    H�\$�=     �
  H�    H�    H�$H�D$   �    H�\$�=     ��  H�    H�    H�$H�D$   �    H�\$�=     �r  H�    H�$    H�    H�\$H�D$   H�    H�\$H�    H�\$ �    H�\$(H�H�$H�KH�L$�    H�\$�=     ��  H�    H�$    H�    H�\$H�D$   H�    H�\$H�    H�\$ �    H�\$(H�H�$H�KH�L$�    H�\$�=     �d  H�    H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     �  H�    1�H��}aH�    H�$H�    H�\$H�    H��Hk�H�H�\$H�    H��H�D$8Hk�H�H�\$H�D$�    H�D$8H��H��|�H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     �?  H�    1�H��}aH�    H�$H�    H�\$H�    H��Hk�H�H�\$H�    H��H�D$8Hk�H�H�\$H�D$�    H�D$8H��H��|�H�    H�$H�D$    H�D$    H�D$    �    H�\$ �=     u|H�    1�H��}aH�    H�$H�    H�\$H�    H��Hk�H�H�\$H�    H��H�D$8Hk�H�H�\$H�D$�    H�D$8H��H��|��    H��@�H�-    H�,$H�\$�    �q���H�-    H�,$H�\$�    ����H�-    H�,$H�\$�    �����H�-    H�,$H�\$�    ����H�-    H�,$H�\$�    ����H�-    H�,$H�\$�    �{���H�-    H�,$H�\$�    �/���H�-    H�,$H�\$�    ������    �8����������̪
      4  "".initdone·   L  "".initdone·   j  "runtime.throwinit   z "".initdone·   �  io.init   �  regexp.init   �  strings.init   �  $text/template.init   �  unicode.init   �  go/ast.init   �  go/token.init   �  path.init   �  strconv.init   �  ""..gostring.1   �  $regexp.MustCompile   � (runtime.writeBarrier   �  "".matchRx   �  0go.string."[^a-zA-Z0-9]"   �  $regexp.MustCompile   � (runtime.writeBarrier   �   "".nonAlphaNumRx   �  Hgo.string."(?i)^[[:space:]]*output:"   �  $regexp.MustCompile   � (runtime.writeBarrier   �  "".outputPrefix   �  (go.string."^[ \\t]*"   �  "".noteMarker   � "".noteMarker   �  *runtime.concatstring2   �  $regexp.MustCompile   � (runtime.writeBarrier   �  "".noteMarkerRx   �  2go.string."^/[/*][ \\t]*"   �  "".noteMarker   � "".noteMarker   �  *runtime.concatstring2   �  $regexp.MustCompile   � (runtime.writeBarrier   �   "".noteCommentRx   �  (type.map[string]bool   �  runtime.makemap   � (runtime.writeBarrier   �  &"".predeclaredTypes   �  (type.map[string]bool   �  &"".predeclaredTypes   �	  """.statictmp_1012   �	  """.statictmp_1012   �	  $runtime.mapassign1   �
  (type.map[string]bool   �
  runtime.makemap   �
 (runtime.writeBarrier   �  &"".predeclaredFuncs   �  (type.map[string]bool   �  &"".predeclaredFuncs   �  """.statictmp_1014   �  """.statictmp_1014   �  $runtime.mapassign1   �  (type.map[string]bool   �  runtime.makemap   � (runtime.writeBarrier   �  ."".predeclaredConstants   �  (type.map[string]bool   �  ."".predeclaredConstants   �  """.statictmp_1016   �  """.statictmp_1016   �  $runtime.mapassign1   � "".initdone·   �  ."".predeclaredConstants   �  .runtime.writebarrierptr   �  &"".predeclaredFuncs   �  .runtime.writebarrierptr   �  &"".predeclaredTypes   �  .runtime.writebarrierptr   �   "".noteCommentRx   �  .runtime.writebarrierptr   �  "".noteMarkerRx   �  .runtime.writebarrierptr   �  "".outputPrefix   �  .runtime.writebarrierptr   �   "".nonAlphaNumRx   �  .runtime.writebarrierptr   �  "".matchRx   �  .runtime.writebarrierptr   �  0runtime.morestack_noctxt    �  "".autotmp_1017  type.int "".autotmp_1015  type.int "".autotmp_1013 type.int (����� 6od2�� ��o-2�2�2�mm�Di&Di@i��!�������O��  4�	 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <$GOROOT/src/go/doc/synopsis.go:$GOROOT/src/go/doc/comment.go:$GOROOT/src/go/doc/example.go8$GOROOT/src/go/doc/reader.go�(type..hash.[8]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_1027 type.int "".autotmp_1026 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[8]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�$type..eq.[8]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1031 ?type.string "".autotmp_1030 type.string "".autotmp_1029 _type.int "".autotmp_1028 Otype.int "".~r2  type.bool "".q type.*[8]string "".p  type.*[8]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�(type..hash.[1]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_1033 type.int "".autotmp_1032 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[1]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�$type..eq.[1]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1037 ?type.string "".autotmp_1036 type.string "".autotmp_1035 _type.int "".autotmp_1034 Otype.int "".~r2  type.bool "".q type.*[1]string "".p  type.*[1]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�2type..hash."".lineWrapper �  �dH�%    H;a�3  H�� H�\$(H�$H�<$ �  H�\$0H�\$�    H�D$H�\$(H�$H�<$ ��   H�$H�D$0H�D$H�D$   �    H�D$H�\$(H�$H�<$ ��   H�$H�D$0H�D$H�D$   �    H�D$H�\$(H�$H�<$ t^H�$ H�D$0H�D$�    H�D$H�\$(H�$H�<$ t,H�$0H�D$0H�D$H�D$   �    H�\$H�\$8H�� É%    �ˉ%    뙉%    �[����%    �����%    ������    ����
      l  "runtime.interhash   �  runtime.memhash   �  runtime.memhash   �  runtime.strhash   �  runtime.memhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  (type.*"".lineWrapper @�?@6?
 � �  5� Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�.type..eq."".lineWrapper �  �dH�%    H;a�v  H��hH�\$xH�� �\  H�H�sH�\$pH�� �?  H�H�SH9��"  H�D$HH�$H�T$PH�T$H�L$XH�L$H�t$`H�t$�    H�T$xH�D$p�\$ �� ��   �X�j@8�tƄ$�    H��h�H�XH�jH9�tƄ$�    H��h�H�p H�H(H��H�R H�C(H9���   H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    H�L$xH�D$p�\$ �� tAH�X0H�i0H9�tƄ$�    H��h�H�X8H�i8H9�tƄ$�    H��h�Ƅ$�   H��h�Ƅ$�    H��h�Ƅ$�    H��hÉ����������    �m����������������
      �  runtime.ifaceeq   �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1041 type.string "".autotmp_1040 _type.string "".autotmp_1039 ?type.io.Writer "".autotmp_1038 type.io.Writer "".~r2  type.bool "".q (type.*"".lineWrapper "".p  (type.*"".lineWrapper h������u����������� � �  s� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·895d0569a38a56443b84805daa09d838   :$GOROOT/src/go/doc/comment.go�$type..hash."".Note �  �dH�%    H;a��   H�� H�\$(H�$H�<$ ��   H�\$0H�\$H�D$   �    H�D$H�\$(H�$H�<$ tUH�$H�D$0H�D$�    H�D$H�\$(H�$H�<$ t#H�$ H�D$0H�D$�    H�\$H�\$8H�� É%    �ԉ%    뢉%    �i����    �4�������

      ~  runtime.memhash   �  runtime.strhash   �  runtime.strhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  type.*"".Note @�?@? � �  >� Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go� type..eq."".Note �  �dH�%    H;a�  H��HH�L$PH�D$XH�H�(H9�t
�D$` H��H�H�YH�hH9�t
�D$` H��H�H�qH�IH�PH�@H9���   H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� t}H�\$PH�� tnH�S H�C(H�\$XH�� tWH�s H�K(H9�u@H�T$(H�$H�D$0H�D$H�t$8H�t$H�L$@H�L$�    �\$ �� t
�D$`H��H��D$` H��HÉ륉��D$` H��H��    ��������
      �   runtime.eqstring   �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1045  type.string "".autotmp_1044  type.string "".autotmp_1043 ?type.string "".autotmp_1042 type.string "".~r2  type.bool "".q type.*"".Note "".p  type.*"".Note D��������	��� � �  �� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�$type..hash."".Func �  �dH�%    H;a�c  H�� H�\$(H�$H�<$ �?  H�\$0H�\$�    H�D$H�\$(H�$H�<$ �  H�$H�D$0H�D$�    H�D$H�\$(H�$H�<$ ��   H�$ H�D$0H�D$H�D$   �    H�D$H�\$(H�$H�<$ ��   H�$(H�D$0H�D$�    H�D$H�\$(H�$H�<$ t^H�$8H�D$0H�D$�    H�D$H�\$(H�$H�<$ t,H�$HH�D$0H�D$H�D$   �    H�\$H�\$8H�� É%    �ˉ%    뙉%    �d����%    �"����%    ������%    �����    ����
      l  runtime.strhash   �  runtime.strhash   �  runtime.memhash   �  runtime.strhash   �  runtime.strhash   �  runtime.memhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  type.*"".Func @�?@B?
 � �  5� Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go� type..eq."".Func �	  �	dH�%    H;a�7  H��HH�\$PH�� �  H�3H�KH�\$XH�� �   H�H�CH9���  H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� ��  H�\$PH�� ��  H�SH�CH�\$XH�� �x  H�sH�KH9��]  H�T$(H�$H�D$0H�D$H�t$8H�t$H�L$@H�L$�    H�L$PH�D$X�\$ �� �  H�Y H�h H9�t
�D$` H��H�H�q(H�I0H�P(H�@0H9���   H�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� ��   H�\$PH�� ��   H�S8H�C@H�\$XH�� txH�s8H�K@H9�uaH�T$(H�$H�D$0H�D$H�t$8H�t$H�L$@H�L$�    �\$ �� t+H�l$PH�]HL�D$XI�hHH9�t
�D$` H��H��D$`H��H��D$` H��HÉ넉�j����D$` H��H��D$` H��HÉ������c����D$` H��HÉ������������    ����������������
      �   runtime.eqstring   �   runtime.eqstring   �   runtime.eqstring   �   runtime.eqstring   �	  0runtime.morestack_noctxt   0�  "".autotmp_1053  type.string "".autotmp_1052  type.string "".autotmp_1051  type.string "".autotmp_1050  type.string "".autotmp_1049  type.string "".autotmp_1048  type.string "".autotmp_1047 ?type.string "".autotmp_1046 type.string "".~r2  type.bool "".q type.*"".Func "".p  type.*"".Func j�������	��	����	����� � �  s� Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�&"".(*methodSet).set  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�\$8H�+H�,$H�\$@H�\$�    H��0��    �X�����������
      x  go.string."doc"   �  *go.string."methodSet"   �  go.string."set"   �  "runtime.panicwrap   �   "".methodSet.set   �  0runtime.morestack_noctxt    `  "".f *type.*go/ast.FuncDecl ""..this  $type.*"".methodSet `�_ � � 
 w9 Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�&"".(*methodSet).add  �	  �	dH�%    H;a�#  H��PH�Y H��tH�|$XH9;uH�#H�\$X1�H9�uEH�    H�$H�D$   H�    H�\$H�D$	   H�    H�\$ H�D$(   �    H�\$XH�+H�D$`H�    H�$H�l$0H�l$H�D$8H�� ��  H�XH�|$H�H�H�KH�O�    H�L$8H�\$ H�1�H9��  H�YHH�hHH9���   1�H9���   H�YHH�hHH9���   H�    H�$�    H�D$H��H�� ��   W�H����    H�\$8H�� ��   H�kH�D$HL�@L�D$H�l$H�-    H�,$�    H�L$8H�D$HH�� tRH�iHH�hHH�D$@H�    H�$H�\$0H�\$H�L$H�|$ tH�D$H�\$@H�\$�    H��PÉ%    �݉ 몉�l���� �J���H�L$@H�    H�$H�\$0H�\$H�L$H�|$ tH�D$H�\$@H�\$�    뢉%    ��� �y����    �����"
      x  go.string."doc"   �  *go.string."methodSet"   �  go.string."add"   �  "runtime.panicwrap   �  "type."".methodSet   �  4runtime.mapaccess1_faststr   �  type."".Func   �  "runtime.newobject   ��  runtime.duffzero   �  type.string   �  (runtime.typedmemmove   �  "type."".methodSet   �  $runtime.mapassign1   �  "type."".methodSet   �  $runtime.mapassign1   �  0runtime.morestack_noctxt    �  "".autotmp_1057  type.*"".Func "".autotmp_1056  type.*"".Func "".autotmp_1055 type.*"".Func "".autotmp_1054 type.*"".Func "".m /type.*"".Func "".mset ?"type."".methodSet "".m type.*"".Func ""..this  $type.*"".methodSet  ����i�
 � �  wO�T} Tgclocals·6412d3717715814cae1af4eeac4eb5d3 Tgclocals·311743cc5ea08f25d41b6a4d25949ffe   <autogenerated>�."".(*exampleByName).Len  �  �dH�%    H;a��   H��0H�Y H��tH�|$8H9;uH�#H�\$81�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$8H�� tH�+H�CH�kH�D$@H��0É���    �T�������
      x  go.string."doc"   �  2go.string."exampleByName"   �  go.string."Len"   �  "runtime.panicwrap   �  0runtime.morestack_noctxt    `  "".~r0 type.int ""..this  ,type.*"".exampleByName `�_`_ � � 
 w9 Tgclocals·3f5c1f818fa7055d0400cecd34057162 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   <autogenerated>�0"".(*exampleByName).Swap  �  �dH�%    H;a�O  H��XH�Y H��tH�|$`H9;uH�#H�\$`1�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$`H�� ��   H�H�KH�kH�l$PH�D$hH�t$pH9���   H��H�+H�l$8H9���   H��H�T$@H�t$0H�L$HH9�siH�,�L�E �=     u9L�H9�s*H��H�l$8�=     uH�+H��X�H�$H�l$�    ���    H�$L�D$�    H�t$0H�T$@H�L$H��    �    �    ��+����    ��������
      x  go.string."doc"   �  2go.string."exampleByName"   �   go.string."Swap"   �  "runtime.panicwrap   � (runtime.writeBarrier   � (runtime.writeBarrier   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  .runtime.writebarrierptr   �  $runtime.panicindex   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   0�  "".autotmp_1059 ? type.*"".Example "".j Otype.int "".s /*type."".exampleByName "".j  type.int "".i type.int ""..this  ,type.*"".exampleByName  ����R� � 
�  w�* Tgclocals·41a13ac73c712c01973b8fe23f62d694 Tgclocals·bade3c5f6d433f8d8fecc50019bf4c85   <autogenerated>�0"".(*exampleByName).Less  �  �dH�%    H;a�
  H��HH�Y H��tH�|$PH9;uH�#H�\$P1�H9�uEH�    H�$H�D$   H�    H�\$H�D$   H�    H�\$ H�D$(   �    H�\$PH�� ��   L�H�SH�kH�l$@H�L$XH�\$`H9�scI�4�H�.H�M H�$H�MH�L$L�L$0H�T$8H9�s5I�4�H�.H�|$H�M H�H�MH�O�    H�\$ H�� ���D$hH��H��    �    ��p����    ��������������
      x  go.string."doc"   �  2go.string."exampleByName"   �   go.string."Less"   �  "runtime.panicwrap   �  "runtime.cmpstring   �  $runtime.panicindex   �  $runtime.panicindex   �  0runtime.morestack_noctxt   @�  
"".s /*type."".exampleByName "".~r2 0type.bool "".j  type.int "".i type.int ""..this  ,type.*"".exampleByName  ����� � �  w� Tgclocals·2fccd208efe70893f9ac8d682812ae72 Tgclocals·790e5cc5051fc0affc980ade09e929ec   <autogenerated>�2type..hash.[2]go/ast.Decl �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  "runtime.interhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_1062 type.int "".autotmp_1061 type.int "".~r2  type.uintptr "".h type.uintptr "".p  (type.*[2]go/ast.Decl PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�.type..eq.[2]go/ast.Decl �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.ifaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_1066 ? type.go/ast.Decl "".autotmp_1065  type.go/ast.Decl "".autotmp_1064 _type.int "".autotmp_1063 Otype.int "".~r2  type.bool "".q (type.*[2]go/ast.Decl "".p  (type.*[2]go/ast.Decl ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�2type..hash.[1]go/ast.Spec �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  "runtime.interhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_1068 type.int "".autotmp_1067 type.int "".~r2  type.uintptr "".h type.uintptr "".p  (type.*[1]go/ast.Spec PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�.type..eq.[1]go/ast.Spec �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$hH�� ��   H��H��H�H�H�sH�\$`H�� tvH��H��H�H�H�SH9�uVH�D$8H�$H�T$@H�T$H�L$HH�L$H�t$PH�t$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �  runtime.ifaceeq   �  0runtime.morestack_noctxt   0�  "".autotmp_1072 ? type.go/ast.Spec "".autotmp_1071  type.go/ast.Spec "".autotmp_1070 _type.int "".autotmp_1069 Otype.int "".~r2  type.bool "".q (type.*[1]go/ast.Spec "".p  (type.*[1]go/ast.Spec ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�(type..hash.[3]string �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��H��H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  runtime.strhash   �  0runtime.morestack_noctxt   0P  
"".autotmp_1074 type.int "".autotmp_1073 type.int "".~r2  type.uintptr "".h type.uintptr "".p  type.*[3]string PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�$type..eq.[3]string �  �dH�%    H;a��   H��X1�H�D$(   H�l$(H9���   H�D$0H�\$`H�� ��   H��H��H�H�3H�KH�\$hH�� tvH��H��H�H�H�CH9�uVH�t$HH�4$H�L$PH�L$H�T$8H�T$H�D$@H�D$�    �\$ �� t H�D$0H��H�l$(H9��n����D$pH��X��D$p H��XÉ놉�c����    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1078 ?type.string "".autotmp_1077 type.string "".autotmp_1076 _type.int "".autotmp_1075 Otype.int "".~r2  type.bool "".q type.*[3]string "".p  type.*[3]string ,����	��� � �  �S Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�Ltype..hash.struct { a string; b bool } �  �dH�%    H;avvH�� H�\$(H�$H�<$ tYH�\$0H�\$�    H�D$H�\$(H�$H�<$ t,H�$H�D$0H�D$H�D$   �    H�\$H�\$8H�� É%    �ˉ%    ��    �q����
      \  runtime.strhash   �  runtime.memhash   �  0runtime.morestack_noctxt   0@  "".~r2  type.uintptr "".h type.uintptr "".p  Btype.*struct { a string; b bool } @_?@? � � 
 -c Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�Htype..eq.struct { a string; b bool } �  �dH�%    H;a��   H��HH�\$PH�� ��   H�3H�KH�\$XH�� txH�H�CH9�ubH�t$8H�4$H�L$@H�L$H�T$(H�T$H�D$0H�D$�    �\$ �� t,H�l$P�]L�D$XA�h@8�t
�D$` H��H��D$`H��H��D$` H��HÉ넉�k����    �;��������������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  
"".autotmp_1080 ?type.string "".autotmp_1079 type.string "".~r2  type.bool "".q Btype.*struct { a string; b bool } "".p  Btype.*struct { a string; b bool } 8����	��	��� � � 
 ke Tgclocals·3bb21ca8fe1d99a3e492463bd711418a Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440   :$GOROOT/src/go/doc/comment.go�Ttype..hash.[20]struct { a string; b bool } �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��Hk�H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  Ltype..hash.struct { a string; b bool }   �  0runtime.morestack_noctxt   0P  
"".autotmp_1082 type.int "".autotmp_1081 type.int "".~r2  type.uintptr "".h type.uintptr "".p  Jtype.*[20]struct { a string; b bool } PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�Ptype..eq.[20]struct { a string; b bool } �  �dH�%    H;a�  H��h1�H�D$(   H�l$(H9���   H�D$0H�L$pH�� ��   H�\$xH��Hk�H�H�� ��   H��Hk�H�H�L$@H�� ��   H�1H�IH�\$8H�� ��   H�H�CH9�uqH�t$XH�4$H�L$`H�L$H�T$HH�T$H�D$PH�D$�    �\$ �� t;H�l$@�]L�D$8A�h@8�u#H�D$0H��H�l$(H9��4���Ƅ$�   H��h�Ƅ$�    H��hÉ�o�����R�����2���������    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1088 ?type.string "".autotmp_1087 type.string "".autotmp_1086 _Btype.*struct { a string; b bool } "".autotmp_1085 OBtype.*struct { a string; b bool } "".autotmp_1084 type.int "".autotmp_1083 otype.int "".~r2  type.bool "".q Jtype.*[20]struct { a string; b bool } "".p  Jtype.*[20]struct { a string; b bool } ,������� � �  �� Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·34eab47d33fa46b254c22cdccfd2dc77   :$GOROOT/src/go/doc/comment.go�Ttype..hash.[15]struct { a string; b bool } �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��Hk�H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  Ltype..hash.struct { a string; b bool }   �  0runtime.morestack_noctxt   0P  
"".autotmp_1090 type.int "".autotmp_1089 type.int "".~r2  type.uintptr "".h type.uintptr "".p  Jtype.*[15]struct { a string; b bool } PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�Ptype..eq.[15]struct { a string; b bool } �  �dH�%    H;a�  H��h1�H�D$(   H�l$(H9���   H�D$0H�L$pH�� ��   H�\$xH��Hk�H�H�� ��   H��Hk�H�H�L$@H�� ��   H�1H�IH�\$8H�� ��   H�H�CH9�uqH�t$XH�4$H�L$`H�L$H�T$HH�T$H�D$PH�D$�    �\$ �� t;H�l$@�]L�D$8A�h@8�u#H�D$0H��H�l$(H9��4���Ƅ$�   H��h�Ƅ$�    H��hÉ�o�����R�����2���������    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1096 ?type.string "".autotmp_1095 type.string "".autotmp_1094 _Btype.*struct { a string; b bool } "".autotmp_1093 OBtype.*struct { a string; b bool } "".autotmp_1092 type.int "".autotmp_1091 otype.int "".~r2  type.bool "".q Jtype.*[15]struct { a string; b bool } "".p  Jtype.*[15]struct { a string; b bool } ,������� � �  �� Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·34eab47d33fa46b254c22cdccfd2dc77   :$GOROOT/src/go/doc/comment.go�Rtype..hash.[4]struct { a string; b bool } �  �dH�%    H;avpH��(H�L$81�H�D$   H�l$H9�}DH�D$ H�\$0H�� t>H��Hk�H�H�$H�L$8H�L$�    H�L$H�D$ H��H�l$H9�|�H�L$@H��(É��    �w����������
      �  Ltype..hash.struct { a string; b bool }   �  0runtime.morestack_noctxt   0P  
"".autotmp_1098 type.int "".autotmp_1097 type.int "".~r2  type.uintptr "".h type.uintptr "".p  Htype.*[4]struct { a string; b bool } PgOPO � � 
 U; Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2 Tgclocals·33cdeccccebe80329f1fdbee7f5874cb   :$GOROOT/src/go/doc/comment.go�Ntype..eq.[4]struct { a string; b bool } �  �dH�%    H;a�  H��h1�H�D$(   H�l$(H9���   H�D$0H�L$pH�� ��   H�\$xH��Hk�H�H�� ��   H��Hk�H�H�L$@H�� ��   H�1H�IH�\$8H�� ��   H�H�CH9�uqH�t$XH�4$H�L$`H�L$H�T$HH�T$H�D$PH�D$�    �\$ �� t;H�l$@�]L�D$8A�h@8�u#H�D$0H��H�l$(H9��4���Ƅ$�   H��h�Ƅ$�    H��hÉ�o�����R�����2���������    ���������
      �   runtime.eqstring   �  0runtime.morestack_noctxt   0�  "".autotmp_1104 ?type.string "".autotmp_1103 type.string "".autotmp_1102 _Btype.*struct { a string; b bool } "".autotmp_1101 OBtype.*struct { a string; b bool } "".autotmp_1100 type.int "".autotmp_1099 otype.int "".~r2  type.bool "".q Htype.*[4]struct { a string; b bool } "".p  Htype.*[4]struct { a string; b bool } ,������� � �  �� Tgclocals·51af24152615272c3d9efc8538f95767 Tgclocals·34eab47d33fa46b254c22cdccfd2dc77   :$GOROOT/src/go/doc/comment.go�Tgclocals·12fc1489b12fcdedb8fc818b7369b5d9              �Tgclocals·13bdb4aeeaf63de3cc223d640262ea59             �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �Tgclocals·88f14b8ca07e3b9e0b9cbc5ca8ee0278 @  @          @   D      E   A    �Tgclocals·2331195bde16ef19bace3004fa98e646 @  @                         �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·b4c25e9b09fd0cf9bb429dcefe91c353             �Tgclocals·6bdcbbfceecc5cba590c8a52e9a888b3 (  (          �       �Tgclocals·cb395d89503762333b1bfb09ba74eb12 (  (                �bgo.string.hdr.",.;:!?+*/=()[]{}_^°&§~%#@<\">\\"                       Zgo.string.",.;:!?+*/=()[]{}_^°&§~%#@<\">\\"   �Zgo.string.",.;:!?+*/=()[]{}_^°&§~%#@<\">\\" @  @,.;:!?+*/=()[]{}_^°&§~%#@<">\  �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·f47057354ec566066f8688a4970cff5a                  �"go.string.hdr."_"                       go.string."_"   �go.string."_"   _  �(go.string.hdr."hdr-"                        go.string."hdr-"   � go.string."hdr-"   
hdr-  �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �Tgclocals·a7d2bdfc04e5cad614b789a6f5ec96df H  H                           �Tgclocals·46ae46c0833abd65a9bd508c0d4723b4 H  H                            �$go.string.hdr."\n"                       go.string."\n"   �go.string."\n"   
  �Tgclocals·f67a1bd37088b83155134772c74a5fc0 �  �   '            �     �     �    �    �    �    �    �    �$   ��    �Tgclocals·3836fb0d9c1e7dd27acd0557fec71b90 h  h                                        �Tgclocals·da53b597af7c02fca1968f95e2ccd079 p  p   (                                         �Tgclocals·a8e198e4544b9f4af27e2179a8f48de0 @  @   	   W   W   W   W   W   W    �Tgclocals·77c75893cdd92181c21e4e3e10e9f609 (  (                 �Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 (  (                �Tgclocals·23e8278e2b69a3a75fa59b23c49ed6ad              �Tgclocals·87d20ce1b58390b294df80b886db78bf             �&go.string.hdr."BUG"                       go.string."BUG"   �go.string."BUG"   BUG  �Tgclocals·b58df2d7616fbb6904d034404c8af93c �  �   *              ʲ      ʲ    � ʲ    � ʲ    � ʲ   @� ʲ   H� ʲ   I� ʲ   I� ʲ   I ʲ   I ʲ   I  ʲ   	  ʲ     ʲ    �Tgclocals·d40f86804c765b65adbc82845c11e455 �  �                                                    �>Jgo.itab.*go/ast.BlockStmt.go/ast.Node     �>@go.itab.*go/ast.File.go/ast.Node     �>Ngo.itab."".exampleByName.sort.Interface     �(go.string.hdr."Test"                        go.string."Test"   � go.string."Test"   
Test  �2go.string.hdr."Benchmark"             	          *go.string."Benchmark"   �*go.string."Benchmark"    Benchmark  �.go.string.hdr."Example"                       &go.string."Example"   �&go.string."Example"   Example  �Tgclocals·57f34913b4e4f52cd021da0277a0692e �  �   &           +�     +�     k�     {�     �      �     } �     m �     -      ) �     1 �     ! �       �       �            �Tgclocals·a0565663444d773a05e50b742a3936f2 �  �                                                       �"go.string.hdr." "                       go.string." "   �go.string." "      �Tgclocals·fad3647538fe088c3f63d28bb4a0e2d7                   �Tgclocals·5cbd57cf8f9b35eac9551b20a42afe1f                  �Tgclocals·709a14768fab2805a378215c02f0d27f              �Tgclocals·1c5a071f4ad97fe89533b360c694a573             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·3260b5c802f633fd6252c227878dd72a                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·6432f8c6a0d23fa7bee6c5d96f21a92a             �>Lgo.itab.*go/ast.ImportSpec.go/ast.Spec     �>Fgo.itab.*go/ast.GenDecl.go/ast.Decl     �>Hgo.itab.*go/ast.FuncDecl.go/ast.Decl     �*go.string.hdr."_test"                       "go.string."_test"   �"go.string."_test"   _test  �"go.string.hdr."."                       go.string."."   �go.string."."   .  �(go.string.hdr."main"                        go.string."main"   � go.string."main"   
main  �Tgclocals·0b5e8d15b1b34de9bb59946bbdd0aacd �  �B   �                                0                                       �                    �                     �                                                                                                                                                                                                                                       �                    �                    �                   `  TUUU   T         `  TUUU   T  @      `  TUUU   T  @@    `  TUUU   T  @@     `  TUUU   D         `  TUUU   D         `  TUUU   D         `  TUUU   D  @@     `  TUUU   D   @ @  `  TUUU   D        `  TUUU   @�        `  TUUU   @ �      	  `  TUUU               `  TUUU   @        `  TUUU   @       	  `  TUUU   @          `  TUUU   @        	  `  TUUU   �        	  `� TUUU   �      	  `� TUUU   �     @	  `� TUUU   �    @	  `� TUUU   ��    	  `� TUUU   �     	  `� TUUU   �       	  `� TUUU   �       	  `� TUUU   �        	  `� TUUU   �        	  `� TUUU   �       	  `� TUUU   �       	  `� TUUU   �      	  `� TUUU   �        	  `  TUUU   �        	 `  TUUU   �          `  TUUU   �         `  TUUU   �          `  TUUU   �          `  TUUU   �@         `  TUUU   �`         `  TUUU   �        `  TUUU   �         `  TUUU   @        `  TUUU    P        `  TUUU    P        a  TUUU    P         a  TUUU             a  TUUU             `  TUUU              `  TUUU    �Tgclocals·ab21a96c86932eb21e674bd4000cfd30 �  �B                                                                                                                                                                                                             �2go.string.hdr."Copyright"             	          *go.string."Copyright"   �*go.string."Copyright"    Copyright  �Tgclocals·6cf11449797bbc22c96eb58e2aa7d4d6 �  �            � ��  �  � �  �    �  � ��  �   �   �  � " �   �      �Tgclocals·93d42c534c9b7817c9d67e4a28433e4e �  �                                                             �Tgclocals·0ce45eb4af445847db003d38f23f3ab0 8  8                   !    �Tgclocals·87c30dc0786889497a80d853dd7fef3f 8  8                      �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·d98f60bd8519d0c68364b2a1d83af357             �Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0 (  (                 �Tgclocals·adb3347b296419e60da36d67f8b7ce43 (  (                �Tgclocals·83ead081cd909acab0dcd88a450c1878                   �Tgclocals·f47057354ec566066f8688a4970cff5a                  �*go.string.hdr."error"                       "go.string."error"   �"go.string."error"   error  �Tgclocals·82a1413d9c726b969ce192c6dcea957e (  (   
              �Tgclocals·37a2283f5c69c342946cad8073b58fca (  (                �Tgclocals·b6cb89307147056cbbf19b02d7f6310a @  @          �   �   �   �   �    �Tgclocals·ba362c851cf6718bcf08a64a3f3a3743 @  @                         �Tgclocals·83ead081cd909acab0dcd88a450c1878                   �Tgclocals·2f2d69f12d345ece4be5273d9b84f0bb                  �Tgclocals·54334d948b35c5006059bc936ec0efb4 @  @          0                �Tgclocals·948a0e540dd9ee4dc893ee9411d99e55 @  @                         �Tgclocals·cb1549917f9fe0533af2fa9f39272c98 x  x           `         	  �	  �	  �	  �  \    %�   �Tgclocals·d696fea639189e6f0ee17af9ebd01687 x  x                                              �>Bgo.itab.*go/ast.Ident.go/ast.Expr     �>Pgo.itab.*go/ast.SelectorExpr.go/ast.Expr     �Tgclocals·e4ca007442f0c3cdda096ebe56a943a8 `  `
   	       �        $                   �Tgclocals·0f0d539f72a0076bd99eb5022e35364d `  `
                                     �Tgclocals·e127204208a449a4bc3afdf4417ef9c1 0  0             2       �Tgclocals·d8668e205667c6ef4f74e27331326ebc 0  0                   �Tgclocals·d3b071704863cbd459bbd46f550e3b94 (  (                 �Tgclocals·f7aa1743939cae014f83a8a2d262049c (  (                �Tgclocals·9d98f0d067a7d5c31416a70b02745cb5 (  (                 �Tgclocals·7e902992778eda5f91d29a3f0c115aee (  (                �Tgclocals·7b90e273048a3c2d112e626ee7e85da5                   �Tgclocals·51af24152615272c3d9efc8538f95767                  �Tgclocals·8fe27e4ff3724ff01c209913c795c44d @  @          �        d       �Tgclocals·bbe2f308595eed0631fb6c42f0ddbda2 @  @                         �Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0 (  (                 �Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc (  (      	   	   	    �Tgclocals·280b01b991f7f5bfaff037b5a4d2aae0 (  (                 �Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc (  (      	   	   	    �Tgclocals·e61e23fa553179df29e88d2b566c0cc1 (  (                 �Tgclocals·0efbc58fefb81b08b9ededd9b41f7cdc (  (      	   	   	    �Tgclocals·6d07ab0a37c299682f1d85b92cb6cfd1      	        �Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6             �"go.string.hdr."*"                       go.string."*"   �go.string."*"   *  �.go.string.hdr."BADRECV"                       &go.string."BADRECV"   �&go.string."BADRECV"   BADRECV  �Tgclocals·bade3c5f6d433f8d8fecc50019bf4c85                   �Tgclocals·aefd16b155593f6f07980a05b297ad1f                  �Tgclocals·c479f047767b723c63a86ea32fdba623 P  P          @   P  P  R         �Tgclocals·cebf12d22eea72c192e5960fe2f61bf0 P  P                               �Tgclocals·008e235a1392cc90d1ed9ad2f7e76d87 (  (                 �Tgclocals·7e902992778eda5f91d29a3f0c115aee (  (                �Tgclocals·21a8f585a14d020f181242c5256583dc                   �Tgclocals·ac82343006770597a842747caad5b201                  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0ebb2d1da58c1b4224bf5a7b370d7578             �Tgclocals·39612780d40568a5b01933408425e52c X  X	   
           0   8   :      
      E    �Tgclocals·573eebd23f15bbede97c85018d63627a X  X	                                  �Tgclocals·e4edfcfe053f06aa2f3f9df5ba415e02 h  h          �   �   �   �   �   �   �   �   	      �Tgclocals·24bdc3afac682cc4abeb732876105abc h  h                                        �Tgclocals·709a14768fab2805a378215c02f0d27f              �Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6             �Tgclocals·0c8aa8e80191a30eac23f1a218103f16                   �Tgclocals·2f2d69f12d345ece4be5273d9b84f0bb                  �Tgclocals·a4ac9012e8051c074b7cac5858bd5519 (  (                �Tgclocals·adb3347b296419e60da36d67f8b7ce43 (  (                �Tgclocals·f76a807c7b8b6a371ade38b5b9694ecd �  �   #           @�      @�                                  %     %     %     %      �                     (                          �Tgclocals·696dc48efaf7c9921882eba1b5b5885e �  �                                                                �Tgclocals·368ff6680f3872f8e014b9f8c1a308ff                   �Tgclocals·f86cabb45f3736e32e1652a4ce443e9b                  �Tgclocals·7301d8fdff8300440e17cffa48be7961 p  p              �  �  �  �  T    !     
    �Tgclocals·e76d9788ffeb8eb69a0d7b2c884b94ed p  p                                           �Tgclocals·e7cc1a3a5ad7e5bd5d4932eddee30345 �  �            	  �	  �	  �	  �  T    !   �     !  �!  �!  �!  �   X      "   �Tgclocals·715f4247ff054ce54b6559cd80f93589 �  �                                                                   �Tgclocals·bddc76d8a57f9840df311eb725104ff2 h  h                 ""   �A !A A   	  �Tgclocals·d40c6564e2ba8bed9102651873b34d14 h  h                                        �Tgclocals·db3311d7e1cb6ec5029186017096a081 (  (                 �Tgclocals·14c16763214c88f6ebc22b4b638329b7 (  (                �>Hgo.itab.*go/ast.TypeSpec.go/ast.Spec     �Tgclocals·3eb79ea418853034459ea0e413208728 �  �   "             `             1       1 �     0       v       ~       ~      >      >       4        �Tgclocals·a21ab7bae19632fedab25371b764faba p  p                                           �Tgclocals·7fe2912721285589731dc5ce1f08c6a7 0  0           �        �Tgclocals·42e7756549fd1f1e78e70fcb9f08dd2b 0  0                   �>Hgo.itab.*go/ast.StarExpr.go/ast.Expr     �Tgclocals·705a498ed8ccdac9185f030fb45a87b7 �  �              $   %   &   "   �  �  �!  �  �  �  �  �  @    �Tgclocals·86c3de611c79526d490a82204ab8e699 �  �                                                    �Tgclocals·ff840c582379ce333f10594801100e10 X  X	                ��?��?��?��?��?� � �Tgclocals·11c63aa4b444ca1a56e95d01623cf60d X  X	      �   �   �   �   �   �   �   �   �    �Tgclocals·81bdb1fcce921ebe87bf14577379b26e P  P   "           ���?    ���?    ��/      �Tgclocals·5d2b5a2aeff4e4cf961f497a12cc05ae 0  0                   �Tgclocals·cf6154774c0aa37b6123d9727e16ac04 �  �   ,               �      �   @ �   H �    ��   ��   # ��    �Tgclocals·a9ea41aae9e32efcc8711d8fabe405fb P  P                               �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �>>go.itab.*"".data.sort.Interface     �Tgclocals·2c033e7f4f4a74cc7e9f368d1fec9f60                   �Tgclocals·51af24152615272c3d9efc8538f95767                  �Tgclocals·ef5fd2c82c386cd66d746b952cc06875 0  0          �  �      �Tgclocals·c87a734079562d73ffd9eee8328c7183 0  0                   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·ad7181e2240ebb348baa41afdc8d0afe 8  8   	             
       �Tgclocals·4a5c83272286258cf484ac950366f973 8  8                      �Tgclocals·748e3f8a785e34acbbe52dd60e6e6e96 �  �           � � � �$��$��$��$��$���� � �  �          �Tgclocals·330a8f52616cf9d268418fab976acddc �  �                                                          �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �Tgclocals·98894f398543f5a4f57ec3edfd994f6a H  H          ��  � �� �   �   �    �Tgclocals·fb63e74b6f2618e7c5d9866e2c2934f2 H  H                            �Tgclocals·3fda2e0c42698195f82d5b8e047ca0ad (  (   	          	    �Tgclocals·adb3347b296419e60da36d67f8b7ce43 (  (                �Tgclocals·d8fdd2a55187867c76648dc792366181                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·89fe65749ce0afc971c0982226501ff0             �Tgclocals·575fdb695a683406ac81277ae7ac66b5 (  (          !       �Tgclocals·55cc6ee7528f0b48e5a6d9bfba36524a (  (                �Tgclocals·9edbfbd6af913bb4812a079f727a5e32 0  0                    �Tgclocals·f6bd6b3389b872033d462029172c8612           �Tgclocals·008e235a1392cc90d1ed9ad2f7e76d87 (  (                 �Tgclocals·9c91d8a91ac42440a3d1507bc8d2e808 (  (                �Tgclocals·ce81e155410342c1a623d0fa5be5f2a2               �    �Tgclocals·f56b2291fa344104975cb6587be42b9b                    �Tgclocals·f304628972275ea37e1ee36ac34113c0                   �Tgclocals·c55cf99de9cdd8c8202a466952fa1a45                    �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·f304628972275ea37e1ee36ac34113c0                   �Tgclocals·c55cf99de9cdd8c8202a466952fa1a45                    �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·f304628972275ea37e1ee36ac34113c0                   �Tgclocals·c55cf99de9cdd8c8202a466952fa1a45                    �>""..gobytes.1   &ldquo; �>""..gobytes.2   &rdquo; �>""..gobytes.3   <a href=" �>""..gobytes.4   "> �>""..gobytes.5   </a> �>""..gobytes.6   <i> �>""..gobytes.7   </i> �>""..gobytes.8   <p>
 �>""..gobytes.9 
  
</p>
 �>""..gobytes.10 
  
<pre> �>""..gobytes.11   </pre>
 �>""..gobytes.12   <h3 id=" �>""..gobytes.13   "> �>""..gobytes.14   </h3>
 �>""..gobytes.15   
 �>""..gobytes.16     �Xgo.string.hdr."([A-Z][A-Z]+)\\(([^)]+)\\):?"                       Pgo.string."([A-Z][A-Z]+)\\(([^)]+)\\):?"   �Pgo.string."([A-Z][A-Z]+)\\(([^)]+)\\):?" @  6([A-Z][A-Z]+)\(([^)]+)\):?  �2go.string.hdr."copyright"             	          *go.string."copyright"   �*go.string."copyright"    copyright  �4go.string.hdr."all rights"             
          ,go.string."all rights"   �,go.string."all rights"    all rights  �,go.string.hdr."author"                       $go.string."author"   �$go.string."author"   author  �$"".hdr..gostring.1             �          ""..gostring.1   �""..gostring.1 �  �((https?|ftp|file|gopher|mailto|news|nntp|telnet|wais|prospero)://[a-zA-Z0-9_@\-]+([.:][a-zA-Z0-9_@\-]+)*/?[a-zA-Z0-9_?%#~&/\-+=()]+([:.,][a-zA-Z0-9_?%#~&/\-+=()]+)*)|([\pL_][\pL_0-9]*)  �8go.string.hdr."[^a-zA-Z0-9]"                       0go.string."[^a-zA-Z0-9]"   �0go.string."[^a-zA-Z0-9]"    [^a-zA-Z0-9]  �Pgo.string.hdr."(?i)^[[:space:]]*output:"                       Hgo.string."(?i)^[[:space:]]*output:"   �Hgo.string."(?i)^[[:space:]]*output:" @  2(?i)^[[:space:]]*output:  �0go.string.hdr."^[ \\t]*"                       (go.string."^[ \\t]*"   �(go.string."^[ \\t]*"   ^[ \t]*  �:go.string.hdr."^/[/*][ \\t]*"                       2go.string."^/[/*][ \\t]*"   �2go.string."^/[/*][ \\t]*"    ^/[/*][ \t]*  �(go.string.hdr."bool"                        go.string."bool"   � go.string."bool"   
bool  �(go.string.hdr."byte"                        go.string."byte"   � go.string."byte"   
byte  �2go.string.hdr."complex64"             	          *go.string."complex64"   �*go.string."complex64"    complex64  �4go.string.hdr."complex128"             
          ,go.string."complex128"   �,go.string."complex128"    complex128  �.go.string.hdr."float32"                       &go.string."float32"   �&go.string."float32"   float32  �.go.string.hdr."float64"                       &go.string."float64"   �&go.string."float64"   float64  �&go.string.hdr."int"                       go.string."int"   �go.string."int"   int  �(go.string.hdr."int8"                        go.string."int8"   � go.string."int8"   
int8  �*go.string.hdr."int16"                       "go.string."int16"   �"go.string."int16"   int16  �*go.string.hdr."int32"                       "go.string."int32"   �"go.string."int32"   int32  �*go.string.hdr."int64"                       "go.string."int64"   �"go.string."int64"   int64  �(go.string.hdr."rune"                        go.string."rune"   � go.string."rune"   
rune  �,go.string.hdr."string"                       $go.string."string"   �$go.string."string"   string  �(go.string.hdr."uint"                        go.string."uint"   � go.string."uint"   
uint  �*go.string.hdr."uint8"                       "go.string."uint8"   �"go.string."uint8"   uint8  �,go.string.hdr."uint16"                       $go.string."uint16"   �$go.string."uint16"   uint16  �,go.string.hdr."uint32"                       $go.string."uint32"   �$go.string."uint32"   uint32  �,go.string.hdr."uint64"                       $go.string."uint64"   �$go.string."uint64"   uint64  �.go.string.hdr."uintptr"                       &go.string."uintptr"   �&go.string."uintptr"   uintptr  �,go.string.hdr."append"                       $go.string."append"   �$go.string."append"   append  �&go.string.hdr."cap"                       go.string."cap"   �go.string."cap"   cap  �*go.string.hdr."close"                       "go.string."close"   �"go.string."close"   close  �.go.string.hdr."complex"                       &go.string."complex"   �&go.string."complex"   complex  �(go.string.hdr."copy"                        go.string."copy"   � go.string."copy"   
copy  �,go.string.hdr."delete"                       $go.string."delete"   �$go.string."delete"   delete  �(go.string.hdr."imag"                        go.string."imag"   � go.string."imag"   
imag  �&go.string.hdr."len"                       go.string."len"   �go.string."len"   len  �(go.string.hdr."make"                        go.string."make"   � go.string."make"   
make  �&go.string.hdr."new"                       go.string."new"   �go.string."new"   new  �*go.string.hdr."panic"                       "go.string."panic"   �"go.string."panic"   panic  �*go.string.hdr."print"                       "go.string."print"   �"go.string."print"   print  �.go.string.hdr."println"                       &go.string."println"   �&go.string."println"   println  �(go.string.hdr."real"                        go.string."real"   � go.string."real"   
real  �.go.string.hdr."recover"                       &go.string."recover"   �&go.string."recover"   recover  �*go.string.hdr."false"                       "go.string."false"   �"go.string."false"   false  �(go.string.hdr."iota"                        go.string."iota"   � go.string."iota"   
iota  �&go.string.hdr."nil"                       go.string."nil"   �go.string."nil"   nil  �(go.string.hdr."true"                        go.string."true"   � go.string."true"   
true  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �:"".ldquo  0type.[]uint8 0                         ""..gobytes.1   �:"".rdquo  0type.[]uint8 0                         ""..gobytes.2   �<"".matchRx  &type.*regexp.Regexp   �:"".html_a  0type.[]uint8 0        	       	          ""..gobytes.3   �:"".html_aq  0type.[]uint8 0                         ""..gobytes.4   �:"".html_enda  0type.[]uint8 0                         ""..gobytes.5   �:"".html_i  0type.[]uint8 0                         ""..gobytes.6   �:"".html_endi  0type.[]uint8 0                         ""..gobytes.7   �:"".html_p  0type.[]uint8 0                         ""..gobytes.8   �:"".html_endp  0type.[]uint8 0                         ""..gobytes.9   �:"".html_pre  0type.[]uint8 0                         ""..gobytes.10   �:"".html_endpre  0type.[]uint8 0                         ""..gobytes.11   �:"".html_h  0type.[]uint8 0                         ""..gobytes.12   �:"".html_hq  0type.[]uint8 0                         ""..gobytes.13   �:"".html_endh  0type.[]uint8 0                         ""..gobytes.14   �< "".nonAlphaNumRx  &type.*regexp.Regexp   �:
"".nl  0type.[]uint8 0                         ""..gobytes.15   �:"".space  0type.[]uint8 0                         ""..gobytes.16   �<"".outputPrefix  &type.*regexp.Regexp   �<"".noteMarker   type.string                    Pgo.string."([A-Z][A-Z]+)\\(([^)]+)\\):?"   �<"".noteMarkerRx  &type.*regexp.Regexp   �< "".noteCommentRx  &type.*regexp.Regexp   �<&"".predeclaredTypes  (type.map[string]bool   �<&"".predeclaredFuncs  (type.map[string]bool   �<."".predeclaredConstants  (type.map[string]bool   �<$"".IllegalPrefixes  0type.[]string 0                         """.statictmp_1011   �<""".statictmp_1011  `type.[3]string `        	               
                         *go.string."copyright"      ,go.string."all rights"   @  $go.string."author"   �>"".initdone·  type.uint8   �""".statictmp_1012  �Htype.[20]struct { a string; b bool } �                                                    	                      
                                                                                                                                                                                                                                                                                                                                                                       (    go.string."bool"   0   go.string."byte"   `  *go.string."complex64"   �  ,go.string."complex128"   �  "go.string."error"   �  &go.string."float32"   �  &go.string."float64"   �  go.string."int"   �   go.string."int8"   �  "go.string."int16"   �  "go.string."int32"   �  "go.string."int64"   �   go.string."rune"   �  $go.string."string"   �   go.string."uint"   �  "go.string."uint8"   �  $go.string."uint16"   �  $go.string."uint32"   �  $go.string."uint64"   �  &go.string."uintptr"   �""".statictmp_1014  �Htype.[15]struct { a string; b bool } �                                                                                                                                                                                                                                                                                                                                      $go.string."append"   0  go.string."cap"   `  "go.string."close"   �  &go.string."complex"   �   go.string."copy"   �  $go.string."delete"   �   go.string."imag"   �  go.string."len"   �   go.string."make"   �  go.string."new"   �  "go.string."panic"   �  "go.string."print"   �  &go.string."println"   �   go.string."real"   �  &go.string."recover"   �""".statictmp_1016  �Ftype.[4]struct { a string; b bool } �                                                                                    "go.string."false"   0   go.string."iota"   `  go.string."nil"   �   go.string."true"   �&"".commentEscape·f               "".commentEscape   �6"".pairedParensPrefixLen·f              0"".pairedParensPrefixLen   �"".emphasize·f              "".emphasize   �"".indentLen·f              "".indentLen   �"".isBlank·f              "".isBlank   �$"".commonPrefix·f              "".commonPrefix   �"".unindent·f              "".unindent   �"".heading·f              "".heading   �"".anchorID·f              "".anchorID   �"".ToHTML·f              "".ToHTML   �"".blocks·f              "".blocks   �"".ToText·f              "".ToText   �4"".(*lineWrapper).write·f              ."".(*lineWrapper).write   �4"".(*lineWrapper).flush·f              ."".(*lineWrapper).flush   �"".New·f              "".New   �"".Examples·f              "".Examples   �&"".exampleOutput·f               "".exampleOutput   �"".isTest·f              "".isTest   �."".exampleByName.Len·f              ("".exampleByName.Len   �0"".exampleByName.Swap·f              *"".exampleByName.Swap   �0"".exampleByName.Less·f              *"".exampleByName.Less   �""".playExample·f              "".playExample   �*"".playExampleFile·f              $"".playExampleFile   �0"".stripOutputComment·f              *"".stripOutputComment   �""".lastComment·f              "".lastComment   �*"".filterIdentList·f              $"".filterIdentList   �*"".hasExportedName·f              $"".hasExportedName   �,"".removeErrorField·f              &"".removeErrorField   �>"".(*reader).filterFieldList·f              8"".(*reader).filterFieldList   �>"".(*reader).filterParamList·f              8"".(*reader).filterParamList   �4"".(*reader).filterType·f              ."".(*reader).filterType   �4"".(*reader).filterSpec·f              ."".(*reader).filterSpec   �&"".copyConstType·f               "".copyConstType   �<"".(*reader).filterSpecList·f              6"".(*reader).filterSpecList   �4"".(*reader).filterDecl·f              ."".(*reader).filterDecl   �6"".(*reader).fileExports·f              0"".(*reader).fileExports   �""".matchFields·f              "".matchFields   �"".matchDecl·f              "".matchDecl   �$"".filterValues·f              "".filterValues   �""".filterFuncs·f              "".filterFuncs   �""".filterTypes·f              "".filterTypes   �."".(*Package).Filter·f              ("".(*Package).Filter   � "".recvString·f              "".recvString   �&"".methodSet.set·f               "".methodSet.set   �&"".methodSet.add·f               "".methodSet.add   �$"".baseTypeName·f              "".baseTypeName   �2"".(*reader).isVisible·f              ,"".(*reader).isVisible   �4"".(*reader).lookupType·f              ."".(*reader).lookupType   �H"".(*reader).recordAnonymousField·f              B"".(*reader).recordAnonymousField   �."".(*reader).readDoc·f              ("".(*reader).readDoc   �0"".(*reader).remember·f              *"".(*reader).remember   �"".specNames·f              "".specNames   �2"".(*reader).readValue·f              ,"".(*reader).readValue   �"".fields·f              "".fields   �0"".(*reader).readType·f              *"".(*reader).readType   �0"".(*reader).readFunc·f              *"".(*reader).readFunc   �0"".(*reader).readNote·f              *"".(*reader).readNote   �2"".(*reader).readNotes·f              ,"".(*reader).readNotes   �0"".(*reader).readFile·f              *"".(*reader).readFile   �6"".(*reader).readPackage·f              0"".(*reader).readPackage   �&"".customizeRecv·f               "".customizeRecv   �L"".(*reader).collectEmbeddedMethods·f              F"".(*reader).collectEmbeddedMethods   �B"".(*reader).computeMethodSets·f              <"".(*reader).computeMethodSets   �8"".(*reader).cleanupTypes·f              2"".(*reader).cleanupTypes   �""".(*data).Len·f              "".(*data).Len   �$"".(*data).Swap·f              "".(*data).Swap   �$"".(*data).Less·f              "".(*data).Less   �"".sortBy·f              "".sortBy   � "".sortedKeys·f              "".sortedKeys   �""".sortingName·f              "".sortingName   �$"".sortedValues·f              "".sortedValues   �""".sortedTypes·f              "".sortedTypes   � "".removeStar·f              "".removeStar   �""".sortedFuncs·f              "".sortedFuncs   � "".noteBodies·f              "".noteBodies   �,"".firstSentenceLen·f              &"".firstSentenceLen   �"".clean·f              "".clean   �"".Synopsis·f              "".Synopsis   �$"".blocks.func1·f              "".blocks.func1   �."".playExample.func1·f              ("".playExample.func1   �0"".sortedValues.func1·f              *"".sortedValues.func1   �0"".sortedValues.func2·f              *"".sortedValues.func2   �."".sortedTypes.func1·f              ("".sortedTypes.func1   �."".sortedTypes.func2·f              ("".sortedTypes.func2   �."".sortedFuncs.func1·f              ("".sortedFuncs.func1   �."".sortedFuncs.func2·f              ("".sortedFuncs.func2   �"".init·f              "".init   �"runtime.gcbits.01    �.go.string.hdr."[]uint8"                       &go.string."[]uint8"   �&go.string."[]uint8"   []uint8  �type.[]uint8 �  �              �~.8                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  .go.string.hdr."[]uint8"   p  *go.weak.type.*[]uint8   �  type.uint8   �6go.typelink.[]uint8	[]uint8              type.[]uint8   �runtime.gcbits.      �0go.string.hdr."[8]uint8"                       (go.string."[8]uint8"   �(go.string."[8]uint8"    [8]uint8  �type.[8]uint8 �  �               >�0� �                                                               0�  runtime.algarray   @  runtime.gcbits.   P  0go.string.hdr."[8]uint8"   p  ,go.weak.type.*[8]uint8   �  type.uint8   �  type.[]uint8   �:go.typelink.[8]uint8	[8]uint8              type.[8]uint8   �0go.string.hdr."[]string"                       (go.string."[]string"   �(go.string."[]string"    []string  �type.[]string �  �              Ө�
                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  0go.string.hdr."[]string"   p  ,go.weak.type.*[]string   �  type.string   �:go.typelink.[]string	[]string              type.[]string   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[8]string              (type..hash.[8]string   �,type..eqfunc.[8]string              $type..eq.[8]string   �&type..alg.[8]string                        0type..hashfunc.[8]string     ,type..eqfunc.[8]string   �&runtime.gcbits.5555   UU �2go.string.hdr."[8]string"             	          *go.string."[8]string"   �*go.string."[8]string"    [8]string  �type.[8]string �  ��       x       US�>                                                                0  &type..alg.[8]string   @  &runtime.gcbits.5555   P  2go.string.hdr."[8]string"   p  .go.weak.type.*[8]string   �  type.string   �  type.[]string   �>go.typelink.[8]string	[8]string              type.[8]string   �Rgo.string.hdr."*map.bucket[string]string"                       Jgo.string."*map.bucket[string]string"   �Jgo.string."*map.bucket[string]string" @  4*map.bucket[string]string  �<type.*map.bucket[string]string �  �              �te 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."*map.bucket[string]string"   p  Ngo.weak.type.**map.bucket[string]string   �  :type.map.bucket[string]string   �2runtime.gcbits.aaaaaaaa02 
  
���� �Pgo.string.hdr."map.bucket[string]string"                       Hgo.string."map.bucket[string]string"   �Hgo.string."map.bucket[string]string" @  2map.bucket[string]string  �.go.string.hdr."topbits"                       &go.string."topbits"   �&go.string."topbits"   topbits  �(go.string.hdr."keys"                        go.string."keys"   � go.string."keys"   
keys  �,go.string.hdr."values"                       $go.string."values"   �$go.string."values"   values  �0go.string.hdr."overflow"                       (go.string."overflow"   �(go.string."overflow"    overflow  �:type.map.bucket[string]string �  �            �>                                                                                                                                                                              �                                             0�  runtime.algarray   @  2runtime.gcbits.aaaaaaaa02   P  Pgo.string.hdr."map.bucket[string]string"   p  Lgo.weak.type.*map.bucket[string]string   �� :type.map.bucket[string]string   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  type.[8]string   �  0go.string.hdr."overflow"   �  <type.*map.bucket[string]string   �"runtime.gcbits.2c   , �Jgo.string.hdr."map.hdr[string]string"                       Bgo.string."map.hdr[string]string"   �Bgo.string."map.hdr[string]string" 0  ,map.hdr[string]string  �*go.string.hdr."count"                       "go.string."count"   �"go.string."count"   count  �*go.string.hdr."flags"                       "go.string."flags"   �"go.string."flags"   flags  �"go.string.hdr."B"                       go.string."B"   �go.string."B"   B  �*go.string.hdr."hash0"                       "go.string."hash0"   �"go.string."hash0"   hash0  �.go.string.hdr."buckets"                       &go.string."buckets"   �&go.string."buckets"   buckets  �4go.string.hdr."oldbuckets"             
          ,go.string."oldbuckets"   �,go.string."oldbuckets"    oldbuckets  �2go.string.hdr."nevacuate"             	          *go.string."nevacuate"   �*go.string."nevacuate"    nevacuate  �4type.map.hdr[string]string �  �0       0       �mlh                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Jgo.string.hdr."map.hdr[string]string"   p  Fgo.weak.type.*map.hdr[string]string   �� 4type.map.hdr[string]string   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  <type.*map.bucket[string]string   �  4go.string.hdr."oldbuckets"   �  <type.*map.bucket[string]string   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �Bgo.string.hdr."map[string]string"                       :go.string."map[string]string"   �:go.string."map[string]string" 0  $map[string]string  �,type.map[string]string �  �              Y��) 5                                                                          0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."map[string]string"   p  >go.weak.type.*map[string]string   �  type.string   �  type.string   �  :type.map.bucket[string]string   �  4type.map.hdr[string]string   �^go.typelink.map[string]string	map[string]string              ,type.map[string]string   �*go.string.hdr."[]int"                       "go.string."[]int"   �"go.string."[]int"   []int  �type.[]int �  �              �f�                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  *go.string.hdr."[]int"   p  &go.weak.type.*[]int   �  type.int   �.go.typelink.[]int	[]int              type.[]int   �.go.string.hdr."*doc.op"                       &go.string."*doc.op"   �&go.string."*doc.op"   *doc.op  �type.*"".op  �  �              �|�� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  .go.string.hdr."*doc.op"   p  (go.weak.type.**"".op   �  type."".op   �,go.string.hdr."doc.op"                       $go.string."doc.op"   �$go.string."doc.op"   doc.op  �$go.string.hdr."op"                       go.string."op"   �go.string."op"   op  �,go.string.hdr."go/doc"                       $go.string."go/doc"   �$go.string."go/doc"   go/doc  �"go.importpath."".                       $go.string."go/doc"   �type."".op  �  �               ��o �                                                                                0�  runtime.algarray   @  runtime.gcbits.   P  ,go.string.hdr."doc.op"   p  type.*"".op   `� type."".op   �  $go.string.hdr."op"   �  "go.importpath."".   �� type."".op   �4go.string.hdr."*doc.block"             
          ,go.string."*doc.block"   �,go.string."*doc.block"    *doc.block  �type.*"".block  �  �              �Ǉ 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*doc.block"   p  .go.weak.type.**"".block   �  type."".block   �"runtime.gcbits.02    �2go.string.hdr."doc.block"             	          *go.string."doc.block"   �*go.string."doc.block"    doc.block  �*go.string.hdr."lines"                       "go.string."lines"   �"go.string."lines"   lines  �*go.string.hdr."block"                       "go.string."block"   �"go.string."block"   block  �type."".block  �  �               @�x                                                                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.02   P  2go.string.hdr."doc.block"   p  type.*"".block   �� type."".block   �  $go.string.hdr."op"   �  "go.importpath."".   �  type."".op   �  *go.string.hdr."lines"   �  "go.importpath."".   �  type.[]string   `� type."".block   �  *go.string.hdr."block"   �  "go.importpath."".   �� type."".block   �6go.string.hdr."[]doc.block"                       .go.string."[]doc.block"   �.go.string."[]doc.block"    []doc.block  �type.[]"".block �  �              `C                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."[]doc.block"   p  0go.weak.type.*[]"".block   �  type."".block   �Dgo.typelink.[]doc.block	[]"".block              type.[]"".block   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �0type..hashfunc.[1]string              (type..hash.[1]string   �,type..eqfunc.[1]string              $type..eq.[1]string   �&type..alg.[1]string                        0type..hashfunc.[1]string     ,type..eqfunc.[1]string   �2go.string.hdr."[1]string"             	          *go.string."[1]string"   �*go.string."[1]string"    [1]string  �type.[1]string �  �              ĸb                                                                 0  &type..alg.[1]string   @  "runtime.gcbits.01   P  2go.string.hdr."[1]string"   p  .go.weak.type.*[1]string   �  type.string   �  type.[]string   �>go.typelink.[1]string	[1]string              type.[1]string   �,go.string.hdr."func()"                       $go.string."func()"   �$go.string."func()"   func()  �type.func() �  �              ���� 3                                                                                                0�  runtime.algarray   @  "runtime.gcbits.01   P  ,go.string.hdr."func()"   p  (go.weak.type.*func()   �� type.func()   �� type.func()   �2go.typelink.func()	func()              type.func()   �2go.string.hdr."*[]string"             	          *go.string."*[]string"   �*go.string."*[]string"    *[]string  �type.*[]string �  �              �"v� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*[]string"   p  .go.weak.type.**[]string   �  type.[]string   �8go.string.hdr."*[]doc.block"                       0go.string."*[]doc.block"   �0go.string."*[]doc.block"    *[]doc.block  � type.*[]"".block �  �              Q� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."*[]doc.block"   p  2go.weak.type.**[]"".block   �  type.[]"".block   � type..hashfunc24                       ,runtime.memhash_varlen   �type..eqfunc24                       .runtime.memequal_varlen   �type..alg24                         type..hashfunc24     type..eqfunc24   �"runtime.gcbits.06    ��go.string.hdr."struct { F uintptr; para *[]string; out *[]doc.block }"             6          �go.string."struct { F uintptr; para *[]string; out *[]doc.block }"   ��go.string."struct { F uintptr; para *[]string; out *[]doc.block }" p  nstruct { F uintptr; para *[]string; out *[]doc.block }  �$go.string.hdr.".F"                       go.string.".F"   �go.string.".F"   .F  �(go.string.hdr."para"                        go.string."para"   � go.string."para"   
para  �&go.string.hdr."out"                       go.string."out"   �go.string."out"   out  �ttype.struct { F uintptr; para *[]string; out *[]"".block } �  �              u^i                                                                                                                                                                                     0  type..alg24   @  "runtime.gcbits.06   P  �go.string.hdr."struct { F uintptr; para *[]string; out *[]doc.block }"   p  �go.weak.type.*struct { F uintptr; para *[]string; out *[]"".block }   �� ttype.struct { F uintptr; para *[]string; out *[]"".block }   �  $go.string.hdr.".F"   �  "go.importpath."".   �  type.uintptr   �  (go.string.hdr."para"   �  "go.importpath."".   �  type.*[]string   �  &go.string.hdr."out"   �  "go.importpath."".   �   type.*[]"".block   ��go.string.hdr."*struct { F uintptr; para *[]string; out *[]doc.block }"             7          �go.string."*struct { F uintptr; para *[]string; out *[]doc.block }"   ��go.string."*struct { F uintptr; para *[]string; out *[]doc.block }" p  p*struct { F uintptr; para *[]string; out *[]doc.block }  �vtype.*struct { F uintptr; para *[]string; out *[]"".block } �  �              ��<0 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."*struct { F uintptr; para *[]string; out *[]doc.block }"   p  �go.weak.type.**struct { F uintptr; para *[]string; out *[]"".block }   �  ttype.struct { F uintptr; para *[]string; out *[]"".block }   �4go.string.hdr."*[1]string"             
          ,go.string."*[1]string"   �,go.string."*[1]string"    *[1]string  �type.*[1]string �  �              l.!� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*[1]string"   p  0go.weak.type.**[1]string   �  type.[1]string   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·895d0569a38a56443b84805daa09d838              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �:type..hashfunc."".lineWrapper              2type..hash."".lineWrapper   �6type..eqfunc."".lineWrapper              .type..eq."".lineWrapper   �0type..alg."".lineWrapper                        :type..hashfunc."".lineWrapper     6type..eqfunc."".lineWrapper   �@go.string.hdr."*doc.lineWrapper"                       8go.string."*doc.lineWrapper"   �8go.string."*doc.lineWrapper" 0  "*doc.lineWrapper  �Lgo.string.hdr."func(*doc.lineWrapper)"                       Dgo.string."func(*doc.lineWrapper)"   �Dgo.string."func(*doc.lineWrapper)" 0  .func(*doc.lineWrapper)  �4type.func(*"".lineWrapper) �  �              L�N 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."func(*doc.lineWrapper)"   p  Fgo.weak.type.*func(*"".lineWrapper)   �� 4type.func(*"".lineWrapper)   �� 4type.func(*"".lineWrapper)   �  (type.*"".lineWrapper   �pgo.typelink.func(*doc.lineWrapper)	func(*"".lineWrapper)              4type.func(*"".lineWrapper)   �\go.string.hdr."func(*doc.lineWrapper, string)"                       Tgo.string."func(*doc.lineWrapper, string)"   �Tgo.string."func(*doc.lineWrapper, string)" @  >func(*doc.lineWrapper, string)  �Dtype.func(*"".lineWrapper, string) �  �              �gr 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(*doc.lineWrapper, string)"   p  Vgo.weak.type.*func(*"".lineWrapper, string)   �� Dtype.func(*"".lineWrapper, string)   �� Dtype.func(*"".lineWrapper, string)   �  (type.*"".lineWrapper   �  type.string   ��go.typelink.func(*doc.lineWrapper, string)	func(*"".lineWrapper, string)              Dtype.func(*"".lineWrapper, string)   �*go.string.hdr."flush"                       "go.string."flush"   �"go.string."flush"   flush  �*go.string.hdr."write"                       "go.string."write"   �"go.string."write"   write  �8go.string.hdr."func(string)"                       0go.string."func(string)"   �0go.string."func(string)"    func(string)  �"type.func(string) �  �              �ǹ� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."func(string)"   p  4go.weak.type.*func(string)   �� "type.func(string)   �� "type.func(string)   �  type.string   �Jgo.typelink.func(string)	func(string)              "type.func(string)   �(type.*"".lineWrapper  �  �              �p}� 6                                                                                                                                                                                      &0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*doc.lineWrapper"   p  :go.weak.type.**"".lineWrapper   �  &type."".lineWrapper   `� (type.*"".lineWrapper   �� (type.*"".lineWrapper   �  *go.string.hdr."flush"   �  "go.importpath."".   �  type.func()   �  4type.func(*"".lineWrapper)   �  ."".(*lineWrapper).flush   �  ."".(*lineWrapper).flush   �  *go.string.hdr."write"   �  "go.importpath."".   �  "type.func(string)   �  Dtype.func(*"".lineWrapper, string)   �  ."".(*lineWrapper).write   �  ."".(*lineWrapper).write   �"runtime.gcbits.13    �>go.string.hdr."doc.lineWrapper"                       6go.string."doc.lineWrapper"   �6go.string."doc.lineWrapper"     doc.lineWrapper  �.go.string.hdr."printed"                       &go.string."printed"   �&go.string."printed"   printed  �*go.string.hdr."width"                       "go.string."width"   �"go.string."width"   width  �,go.string.hdr."indent"                       $go.string."indent"   �$go.string."indent"   indent  �"go.string.hdr."n"                       go.string."n"   �go.string."n"   n  �2go.string.hdr."pendSpace"             	          *go.string."pendSpace"   �*go.string."pendSpace"    pendSpace  �6go.string.hdr."lineWrapper"                       .go.string."lineWrapper"   �.go.string."lineWrapper"    lineWrapper  �&type."".lineWrapper  �  �@       (       2dT%                                                                                                                                                                                                                                                             0                                       8                                               60  0type..alg."".lineWrapper   @  "runtime.gcbits.13   P  >go.string.hdr."doc.lineWrapper"   p  (type.*"".lineWrapper   �� &type."".lineWrapper   �  &go.string.hdr."out"   �  "go.importpath."".   �  type.io.Writer   �  .go.string.hdr."printed"   �  "go.importpath."".   �  type.bool   �  *go.string.hdr."width"   �  "go.importpath."".   �  type.int   �  ,go.string.hdr."indent"   �  "go.importpath."".   �  type.string   �  "go.string.hdr."n"   �  "go.importpath."".   �  type.int   �  2go.string.hdr."pendSpace"   �  "go.importpath."".   �  type.int   `� &type."".lineWrapper   �  6go.string.hdr."lineWrapper"   �  "go.importpath."".   �� &type."".lineWrapper   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �,type..hashfunc."".Note              $type..hash."".Note   �(type..eqfunc."".Note               type..eq."".Note   �"type..alg."".Note                        ,type..hashfunc."".Note     (type..eqfunc."".Note   �"runtime.gcbits.14    �0go.string.hdr."doc.Note"                       (go.string."doc.Note"   �(go.string."doc.Note"    doc.Note  �&go.string.hdr."Pos"                       go.string."Pos"   �go.string."Pos"   Pos  �&go.string.hdr."End"                       go.string."End"   �go.string."End"   End  �&go.string.hdr."UID"                       go.string."UID"   �go.string."UID"   UID  �(go.string.hdr."Body"                        go.string."Body"   � go.string."Body"   
Body  �(go.string.hdr."Note"                        go.string."Note"   � go.string."Note"   
Note  �type."".Note  �  �0       (       �%3                                                                                                                                                                                                                                                                     "0  "type..alg."".Note   @  "runtime.gcbits.14   P  0go.string.hdr."doc.Note"   p  type.*"".Note   �� type."".Note   �  &go.string.hdr."Pos"   �  "type.go/token.Pos   �  &go.string.hdr."End"   �  "type.go/token.Pos   �  &go.string.hdr."UID"   �  type.string   �  (go.string.hdr."Body"   �  type.string   `� type."".Note   �  (go.string.hdr."Note"   �  "go.importpath."".   �� type."".Note   �2go.string.hdr."*doc.Note"             	          *go.string."*doc.Note"   �*go.string."*doc.Note"    *doc.Note  �type.*"".Note  �  �              ��� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*doc.Note"   p  ,go.weak.type.**"".Note   �  type."".Note   �6go.string.hdr."[]*doc.Note"                       .go.string."[]*doc.Note"   �.go.string."[]*doc.Note"    []*doc.Note  �type.[]*"".Note �  �              ��
z                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."[]*doc.Note"   p  0go.weak.type.*[]*"".Note   �  type.*"".Note   �Dgo.typelink.[]*doc.Note	[]*"".Note              type.[]*"".Note   �:go.string.hdr."[][]*doc.Note"                       2go.string."[][]*doc.Note"   �2go.string."[][]*doc.Note"    [][]*doc.Note  �"type.[][]*"".Note �  �              �+                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."[][]*doc.Note"   p  4go.weak.type.*[][]*"".Note   �  type.[]*"".Note   �Lgo.typelink.[][]*doc.Note	[][]*"".Note              "type.[][]*"".Note   �*runtime.gcbits.499224   I�$ �<go.string.hdr."[8][]*doc.Note"                       4go.string."[8][]*doc.Note"   �4go.string."[8][]*doc.Note"    [8][]*doc.Note  �$type.[8][]*"".Note �  ��       �       `2H                                                                0�  runtime.algarray   @  *runtime.gcbits.499224   P  <go.string.hdr."[8][]*doc.Note"   p  6go.weak.type.*[8][]*"".Note   �  type.[]*"".Note   �  "type.[][]*"".Note   �Pgo.typelink.[8][]*doc.Note	[8][]*"".Note              $type.[8][]*"".Note   �\go.string.hdr."*map.bucket[string][]*doc.Note"                       Tgo.string."*map.bucket[string][]*doc.Note"   �Tgo.string."*map.bucket[string][]*doc.Note" @  >*map.bucket[string][]*doc.Note  �Dtype.*map.bucket[string][]*"".Note �  �              � 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."*map.bucket[string][]*doc.Note"   p  Vgo.weak.type.**map.bucket[string][]*"".Note   �  Btype.map.bucket[string][]*"".Note   �6runtime.gcbits.aaaa92244902   ���$I �Zgo.string.hdr."map.bucket[string][]*doc.Note"                       Rgo.string."map.bucket[string][]*doc.Note"   �Rgo.string."map.bucket[string][]*doc.Note" @  <map.bucket[string][]*doc.Note  �Btype.map.bucket[string][]*"".Note �  �P      P      ^���                                                                                                                                                                              �                                       H      0�  runtime.algarray   @  6runtime.gcbits.aaaa92244902   P  Zgo.string.hdr."map.bucket[string][]*doc.Note"   p  Tgo.weak.type.*map.bucket[string][]*"".Note   �� Btype.map.bucket[string][]*"".Note   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  $type.[8][]*"".Note   �  0go.string.hdr."overflow"   �  Dtype.*map.bucket[string][]*"".Note   �Tgo.string.hdr."map.hdr[string][]*doc.Note"                       Lgo.string."map.hdr[string][]*doc.Note"   �Lgo.string."map.hdr[string][]*doc.Note" @  6map.hdr[string][]*doc.Note  �<type.map.hdr[string][]*"".Note �  �0       0       ��                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Tgo.string.hdr."map.hdr[string][]*doc.Note"   p  Ngo.weak.type.*map.hdr[string][]*"".Note   �� <type.map.hdr[string][]*"".Note   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  Dtype.*map.bucket[string][]*"".Note   �  4go.string.hdr."oldbuckets"   �  Dtype.*map.bucket[string][]*"".Note   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �Lgo.string.hdr."map[string][]*doc.Note"                       Dgo.string."map[string][]*doc.Note"   �Dgo.string."map[string][]*doc.Note" 0  .map[string][]*doc.Note  �4type.map[string][]*"".Note �  �              -=� 5                                                                          P0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."map[string][]*doc.Note"   p  Fgo.weak.type.*map[string][]*"".Note   �  type.string   �  type.[]*"".Note   �  Btype.map.bucket[string][]*"".Note   �  <type.map.hdr[string][]*"".Note   �pgo.typelink.map[string][]*doc.Note	map[string][]*"".Note              4type.map[string][]*"".Note   �"runtime.gcbits.25   % �2go.string.hdr."doc.Value"             	          *go.string."doc.Value"   �*go.string."doc.Value"    doc.Value  �&go.string.hdr."Doc"                       go.string."Doc"   �go.string."Doc"   Doc  �*go.string.hdr."Names"                       "go.string."Names"   �"go.string."Names"   Names  �(go.string.hdr."Decl"                        go.string."Decl"   � go.string."Decl"   
Decl  �*go.string.hdr."order"                       "go.string."order"   �"go.string."order"   order  �*go.string.hdr."Value"                       "go.string."Value"   �"go.string."Value"   Value  �type."".Value  �  �8       0       �                                                                                                                                                                              (                                       0                                               $0�  runtime.algarray   @  "runtime.gcbits.25   P  2go.string.hdr."doc.Value"   p  type.*"".Value   �� type."".Value   �  &go.string.hdr."Doc"   �  type.string   �  *go.string.hdr."Names"   �  type.[]string   �  (go.string.hdr."Decl"   �  (type.*go/ast.GenDecl   �  *go.string.hdr."order"   �  "go.importpath."".   �  type.int   `� type."".Value   �  *go.string.hdr."Value"   �  "go.importpath."".   �� type."".Value   �4go.string.hdr."*doc.Value"             
          ,go.string."*doc.Value"   �,go.string."*doc.Value"    *doc.Value  �type.*"".Value  �  �              ��� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."*doc.Value"   p  .go.weak.type.**"".Value   �  type."".Value   �8go.string.hdr."[]*doc.Value"                       0go.string."[]*doc.Value"   �0go.string."[]*doc.Value"    []*doc.Value  � type.[]*"".Value �  �              �0P�                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."[]*doc.Value"   p  2go.weak.type.*[]*"".Value   �  type.*"".Value   �Hgo.typelink.[]*doc.Value	[]*"".Value               type.[]*"".Value   �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·0b86ef39f3fed835f14ba5f4d7c62fa2             �Tgclocals·a8eabfc4a4514ed6b3b0c61e9680e440              �Tgclocals·3bb21ca8fe1d99a3e492463bd711418a             �,type..hashfunc."".Func              $type..hash."".Func   �(type..eqfunc."".Func               type..eq."".Func   �"type..alg."".Func                        ,type..hashfunc."".Func     (type..eqfunc."".Func   �"runtime.gcbits.b5   � �0go.string.hdr."doc.Func"                       (go.string."doc.Func"   �(go.string."doc.Func"    doc.Func  �(go.string.hdr."Name"                        go.string."Name"   � go.string."Name"   
Name  �(go.string.hdr."Recv"                        go.string."Recv"   � go.string."Recv"   
Recv  �(go.string.hdr."Orig"                        go.string."Orig"   � go.string."Orig"   
Orig  �*go.string.hdr."Level"                       "go.string."Level"   �"go.string."Level"   Level  �(go.string.hdr."Func"                        go.string."Func"   � go.string."Func"   
Func  �type."".Func  �  �P       @       �n�                                                                                                                                                                                                                      (                                       8                                       H                                               *0  "type..alg."".Func   @  "runtime.gcbits.b5   P  0go.string.hdr."doc.Func"   p  type.*"".Func   �� type."".Func   �  &go.string.hdr."Doc"   �  type.string   �  (go.string.hdr."Name"   �  type.string   �  (go.string.hdr."Decl"   �  *type.*go/ast.FuncDecl   �  (go.string.hdr."Recv"   �  type.string   �  (go.string.hdr."Orig"   �  type.string   �  *go.string.hdr."Level"   �  type.int   `� type."".Func   �  (go.string.hdr."Func"   �  "go.importpath."".   �� type."".Func   �2go.string.hdr."*doc.Func"             	          *go.string."*doc.Func"   �*go.string."*doc.Func"    *doc.Func  �type.*"".Func  �  �              ܉�� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*doc.Func"   p  ,go.weak.type.**"".Func   �  type."".Func   �6go.string.hdr."[]*doc.Func"                       .go.string."[]*doc.Func"   �.go.string."[]*doc.Func"    []*doc.Func  �type.[]*"".Func �  �              �Q                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."[]*doc.Func"   p  0go.weak.type.*[]*"".Func   �  type.*"".Func   �Dgo.typelink.[]*doc.Func	[]*"".Func              type.[]*"".Func   �&runtime.gcbits.3549   5I �0go.string.hdr."doc.Type"                       (go.string."doc.Type"   �(go.string."doc.Type"    doc.Type  �,go.string.hdr."Consts"                       $go.string."Consts"   �$go.string."Consts"   Consts  �(go.string.hdr."Vars"                        go.string."Vars"   � go.string."Vars"   
Vars  �*go.string.hdr."Funcs"                       "go.string."Funcs"   �"go.string."Funcs"   Funcs  �.go.string.hdr."Methods"                       &go.string."Methods"   �&go.string."Methods"   Methods  �(go.string.hdr."Type"                        go.string."Type"   � go.string."Type"   
Type  �type."".Type  �  ��       x       �h��                                                                                                                                                                                                                      (                                       @                                       X                                       p                                               .0�  runtime.algarray   @  &runtime.gcbits.3549   P  0go.string.hdr."doc.Type"   p  type.*"".Type   �� type."".Type   �  &go.string.hdr."Doc"   �  type.string   �  (go.string.hdr."Name"   �  type.string   �  (go.string.hdr."Decl"   �  (type.*go/ast.GenDecl   �  ,go.string.hdr."Consts"   �   type.[]*"".Value   �  (go.string.hdr."Vars"   �   type.[]*"".Value   �  *go.string.hdr."Funcs"   �  type.[]*"".Func   �  .go.string.hdr."Methods"   �  type.[]*"".Func   `� type."".Type   �  (go.string.hdr."Type"   �  "go.importpath."".   �� type."".Type   �2go.string.hdr."*doc.Type"             	          *go.string."*doc.Type"   �*go.string."*doc.Type"    *doc.Type  �type.*"".Type  �  �              z�Ne 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*doc.Type"   p  ,go.weak.type.**"".Type   �  type."".Type   �6go.string.hdr."[]*doc.Type"                       .go.string."[]*doc.Type"   �.go.string."[]*doc.Type"    []*doc.Type  �type.[]*"".Type �  �              '�t                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."[]*doc.Type"   p  0go.weak.type.*[]*"".Type   �  type.*"".Type   �Dgo.typelink.[]*doc.Type	[]*"".Type              type.[]*"".Type   �8go.string.hdr."*doc.Package"                       0go.string."*doc.Package"   �0go.string."*doc.Package"    *doc.Package  �6go.string.hdr."*doc.Filter"                       .go.string."*doc.Filter"   �.go.string."*doc.Filter"    *doc.Filter  �type.*"".Filter  �  �              ��	q 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."*doc.Filter"   p  0go.weak.type.**"".Filter   �  type."".Filter   �4go.string.hdr."doc.Filter"             
          ,go.string."doc.Filter"   �,go.string."doc.Filter"    doc.Filter  �,go.string.hdr."Filter"                       $go.string."Filter"   �$go.string."Filter"   Filter  �type."".Filter  �  �              g�o 3                                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."doc.Filter"   p  type.*"".Filter   �� type."".Filter   �� type."".Filter   �  type.string   �  type.bool   `� type."".Filter   �  ,go.string.hdr."Filter"   �  "go.importpath."".   �� type."".Filter   �\go.string.hdr."func(*doc.Package, doc.Filter)"                       Tgo.string."func(*doc.Package, doc.Filter)"   �Tgo.string."func(*doc.Package, doc.Filter)" @  >func(*doc.Package, doc.Filter)  �Btype.func(*"".Package, "".Filter) �  �              A��� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(*doc.Package, doc.Filter)"   p  Tgo.weak.type.*func(*"".Package, "".Filter)   �� Btype.func(*"".Package, "".Filter)   �� Btype.func(*"".Package, "".Filter)   �   type.*"".Package   �  type."".Filter   ��go.typelink.func(*doc.Package, doc.Filter)	func(*"".Package, "".Filter)              Btype.func(*"".Package, "".Filter)   �@go.string.hdr."func(doc.Filter)"                       8go.string."func(doc.Filter)"   �8go.string."func(doc.Filter)" 0  "func(doc.Filter)  �(type.func("".Filter) �  �              �=� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."func(doc.Filter)"   p  :go.weak.type.*func("".Filter)   �� (type.func("".Filter)   �� (type.func("".Filter)   �  type."".Filter   �Xgo.typelink.func(doc.Filter)	func("".Filter)              (type.func("".Filter)   � type.*"".Package  �  �              ١z� 6                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."*doc.Package"   p  2go.weak.type.**"".Package   �  type."".Package   `�  type.*"".Package   ��  type.*"".Package   �  ,go.string.hdr."Filter"   �  (type.func("".Filter)   �  Btype.func(*"".Package, "".Filter)   �  ("".(*Package).Filter   �  ("".(*Package).Filter   �.runtime.gcbits.55324902   U2I �6go.string.hdr."doc.Package"                       .go.string."doc.Package"   �.go.string."doc.Package"    doc.Package  �4go.string.hdr."ImportPath"             
          ,go.string."ImportPath"   �,go.string."ImportPath"    ImportPath  �.go.string.hdr."Imports"                       &go.string."Imports"   �&go.string."Imports"   Imports  �2go.string.hdr."Filenames"             	          *go.string."Filenames"   �*go.string."Filenames"    Filenames  �*go.string.hdr."Notes"                       "go.string."Notes"   �"go.string."Notes"   Notes  �(go.string.hdr."Bugs"                        go.string."Bugs"   � go.string."Bugs"   
Bugs  �*go.string.hdr."Types"                       "go.string."Types"   �"go.string."Types"   Types  �.go.string.hdr."Package"                       &go.string."Package"   �&go.string."Package"   Package  �type."".Package  �  ��       �       �8VM                                                                                                                                                                                                                      0                                       H                                       `                                       h                                       �                                       �                                       �                                       �                                               >0�  runtime.algarray   @  .runtime.gcbits.55324902   P  6go.string.hdr."doc.Package"   p   type.*"".Package   �� type."".Package   �  &go.string.hdr."Doc"   �  type.string   �  (go.string.hdr."Name"   �  type.string   �  4go.string.hdr."ImportPath"   �  type.string   �  .go.string.hdr."Imports"   �  type.[]string   �  2go.string.hdr."Filenames"   �  type.[]string   �  *go.string.hdr."Notes"   �  4type.map[string][]*"".Note   �  (go.string.hdr."Bugs"   �  type.[]string   �  ,go.string.hdr."Consts"   �   type.[]*"".Value   �  *go.string.hdr."Types"   �  type.[]*"".Type   �  (go.string.hdr."Vars"   �   type.[]*"".Value   �  *go.string.hdr."Funcs"   �  type.[]*"".Func   `� type."".Package   �  .go.string.hdr."Package"   �  "go.importpath."".   �� type."".Package   �2go.string.hdr."*doc.Mode"             	          *go.string."*doc.Mode"   �*go.string."*doc.Mode"    *doc.Mode  �type.*"".Mode  �  �              ��K 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  2go.string.hdr."*doc.Mode"   p  ,go.weak.type.**"".Mode   �  type."".Mode   �0go.string.hdr."doc.Mode"                       (go.string."doc.Mode"   �(go.string."doc.Mode"    doc.Mode  �(go.string.hdr."Mode"                        go.string."Mode"   � go.string."Mode"   
Mode  �type."".Mode  �  �               ��Y �                                                                                0�  runtime.algarray   @  runtime.gcbits.   P  0go.string.hdr."doc.Mode"   p  type.*"".Mode   `� type."".Mode   �  (go.string.hdr."Mode"   �  "go.importpath."".   �� type."".Mode   � type..hashfunc64             @          ,runtime.memhash_varlen   �type..eqfunc64             @          .runtime.memequal_varlen   �type..alg64                         type..hashfunc64     type..eqfunc64   �,go.string.hdr."[8]int"                       $go.string."[8]int"   �$go.string."[8]int"   [8]int  �type.[8]int �  �@               ��� �                                                               0  type..alg64   @  runtime.gcbits.   P  ,go.string.hdr."[8]int"   p  (go.weak.type.*[8]int   �  type.int   �  type.[]int   �2go.typelink.[8]int	[8]int              type.[8]int   �Lgo.string.hdr."*map.bucket[string]int"                       Dgo.string."*map.bucket[string]int"   �Dgo.string."*map.bucket[string]int" 0  .*map.bucket[string]int  �6type.*map.bucket[string]int �  �              ɾ̜ 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Lgo.string.hdr."*map.bucket[string]int"   p  Hgo.weak.type.**map.bucket[string]int   �  4type.map.bucket[string]int   �.runtime.gcbits.aaaa0002   ��  �Jgo.string.hdr."map.bucket[string]int"                       Bgo.string."map.bucket[string]int"   �Bgo.string."map.bucket[string]int" 0  ,map.bucket[string]int  �4type.map.bucket[string]int �  ��       �       ]hcq                                                                                                                                                                              �                                       �       0�  runtime.algarray   @  .runtime.gcbits.aaaa0002   P  Jgo.string.hdr."map.bucket[string]int"   p  Fgo.weak.type.*map.bucket[string]int   �� 4type.map.bucket[string]int   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  type.[8]int   �  0go.string.hdr."overflow"   �  6type.*map.bucket[string]int   �Dgo.string.hdr."map.hdr[string]int"                       <go.string."map.hdr[string]int"   �<go.string."map.hdr[string]int" 0  &map.hdr[string]int  �.type.map.hdr[string]int �  �0       0       5F�                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Dgo.string.hdr."map.hdr[string]int"   p  @go.weak.type.*map.hdr[string]int   �� .type.map.hdr[string]int   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  6type.*map.bucket[string]int   �  4go.string.hdr."oldbuckets"   �  6type.*map.bucket[string]int   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �<go.string.hdr."map[string]int"                       4go.string."map[string]int"   �4go.string."map[string]int"    map[string]int  �&type.map[string]int �  �              ���J 5                                                                          � 0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."map[string]int"   p  8go.weak.type.*map[string]int   �  type.string   �  type.int   �  4type.map.bucket[string]int   �  .type.map.hdr[string]int   �Rgo.typelink.map[string]int	map[string]int              &type.map[string]int   �@go.string.hdr."[]*doc.namedType"                       8go.string."[]*doc.namedType"   �8go.string."[]*doc.namedType" 0  "[]*doc.namedType  �(type.[]*"".namedType �  �              Pђa                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."[]*doc.namedType"   p  :go.weak.type.*[]*"".namedType   �  $type.*"".namedType   �Xgo.typelink.[]*doc.namedType	[]*"".namedType              (type.[]*"".namedType   �"runtime.gcbits.ff   � �Bgo.string.hdr."[8]*doc.namedType"                       :go.string."[8]*doc.namedType"   �:go.string."[8]*doc.namedType" 0  $[8]*doc.namedType  �*type.[8]*"".namedType �  �@       @       �0�                                                                0  type..alg64   @  "runtime.gcbits.ff   P  Bgo.string.hdr."[8]*doc.namedType"   p  <go.weak.type.*[8]*"".namedType   �  $type.*"".namedType   �  (type.[]*"".namedType   �\go.typelink.[8]*doc.namedType	[8]*"".namedType              *type.[8]*"".namedType   �,go.string.hdr."[]bool"                       $go.string."[]bool"   �$go.string."[]bool"   []bool  �type.[]bool �  �              ���                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  ,go.string.hdr."[]bool"   p  (go.weak.type.*[]bool   �  type.bool   �2go.typelink.[]bool	[]bool              type.[]bool   �.go.string.hdr."[8]bool"                       &go.string."[8]bool"   �&go.string."[8]bool"   [8]bool  �type.[8]bool �  �               s�5 �                                                               0�  runtime.algarray   @  runtime.gcbits.   P  .go.string.hdr."[8]bool"   p  *go.weak.type.*[8]bool   �  type.bool   �  type.[]bool   �6go.typelink.[8]bool	[8]bool              type.[8]bool   �^go.string.hdr."*map.bucket[*doc.namedType]bool"                       Vgo.string."*map.bucket[*doc.namedType]bool"   �Vgo.string."*map.bucket[*doc.namedType]bool" @  @*map.bucket[*doc.namedType]bool  �Ftype.*map.bucket[*"".namedType]bool �  �              e^� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."*map.bucket[*doc.namedType]bool"   p  Xgo.weak.type.**map.bucket[*"".namedType]bool   �  Dtype.map.bucket[*"".namedType]bool   �&runtime.gcbits.fe05   � �\go.string.hdr."map.bucket[*doc.namedType]bool"                       Tgo.string."map.bucket[*doc.namedType]bool"   �Tgo.string."map.bucket[*doc.namedType]bool" @  >map.bucket[*doc.namedType]bool  �Dtype.map.bucket[*"".namedType]bool �  �X       X       ��                                                                                                                                                                              H                                       P       0�  runtime.algarray   @  &runtime.gcbits.fe05   P  \go.string.hdr."map.bucket[*doc.namedType]bool"   p  Vgo.weak.type.*map.bucket[*"".namedType]bool   �� Dtype.map.bucket[*"".namedType]bool   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  *type.[8]*"".namedType   �  ,go.string.hdr."values"   �  type.[8]bool   �  0go.string.hdr."overflow"   �  Ftype.*map.bucket[*"".namedType]bool   �Vgo.string.hdr."map.hdr[*doc.namedType]bool"                       Ngo.string."map.hdr[*doc.namedType]bool"   �Ngo.string."map.hdr[*doc.namedType]bool" @  8map.hdr[*doc.namedType]bool  �>type.map.hdr[*"".namedType]bool �  �0       0       � ��                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Vgo.string.hdr."map.hdr[*doc.namedType]bool"   p  Pgo.weak.type.*map.hdr[*"".namedType]bool   �� >type.map.hdr[*"".namedType]bool   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  Ftype.*map.bucket[*"".namedType]bool   �  4go.string.hdr."oldbuckets"   �  Ftype.*map.bucket[*"".namedType]bool   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �@go.string.hdr."*doc.embeddedSet"                       8go.string."*doc.embeddedSet"   �8go.string."*doc.embeddedSet" 0  "*doc.embeddedSet  �(type.*"".embeddedSet  �  �              �A� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  @go.string.hdr."*doc.embeddedSet"   p  :go.weak.type.**"".embeddedSet   �  &type."".embeddedSet   �>go.string.hdr."doc.embeddedSet"                       6go.string."doc.embeddedSet"   �6go.string."doc.embeddedSet"     doc.embeddedSet  �6go.string.hdr."embeddedSet"                       .go.string."embeddedSet"   �.go.string."embeddedSet"    embeddedSet  �&type."".embeddedSet  �  �              � 5                                                                          X                                          0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."doc.embeddedSet"   p  (type.*"".embeddedSet   �  $type.*"".namedType   �  type.bool   �  Dtype.map.bucket[*"".namedType]bool   �  >type.map.hdr[*"".namedType]bool   `� &type."".embeddedSet   �  6go.string.hdr."embeddedSet"   �  "go.importpath."".   �� &type."".embeddedSet   �8go.string.hdr."[8]*doc.Func"                       0go.string."[8]*doc.Func"   �0go.string."[8]*doc.Func"    [8]*doc.Func  � type.[8]*"".Func �  �@       @       �LLJ                                                                0  type..alg64   @  "runtime.gcbits.ff   P  8go.string.hdr."[8]*doc.Func"   p  2go.weak.type.*[8]*"".Func   �  type.*"".Func   �  type.[]*"".Func   �Hgo.typelink.[8]*doc.Func	[8]*"".Func               type.[8]*"".Func   �Xgo.string.hdr."*map.bucket[string]*doc.Func"                       Pgo.string."*map.bucket[string]*doc.Func"   �Pgo.string."*map.bucket[string]*doc.Func" @  :*map.bucket[string]*doc.Func  �@type.*map.bucket[string]*"".Func �  �              �
�� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."*map.bucket[string]*doc.Func"   p  Rgo.weak.type.**map.bucket[string]*"".Func   �  >type.map.bucket[string]*"".Func   �.runtime.gcbits.aaaafe03   ��� �Vgo.string.hdr."map.bucket[string]*doc.Func"                       Ngo.string."map.bucket[string]*doc.Func"   �Ngo.string."map.bucket[string]*doc.Func" @  8map.bucket[string]*doc.Func  �>type.map.bucket[string]*"".Func �  ��       �       �H�                                                                                                                                                                              �                                       �       0�  runtime.algarray   @  .runtime.gcbits.aaaafe03   P  Vgo.string.hdr."map.bucket[string]*doc.Func"   p  Pgo.weak.type.*map.bucket[string]*"".Func   �� >type.map.bucket[string]*"".Func   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �   type.[8]*"".Func   �  0go.string.hdr."overflow"   �  @type.*map.bucket[string]*"".Func   �Pgo.string.hdr."map.hdr[string]*doc.Func"                       Hgo.string."map.hdr[string]*doc.Func"   �Hgo.string."map.hdr[string]*doc.Func" @  2map.hdr[string]*doc.Func  �8type.map.hdr[string]*"".Func �  �0       0       �[�K                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Pgo.string.hdr."map.hdr[string]*doc.Func"   p  Jgo.weak.type.*map.hdr[string]*"".Func   �� 8type.map.hdr[string]*"".Func   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  @type.*map.bucket[string]*"".Func   �  4go.string.hdr."oldbuckets"   �  @type.*map.bucket[string]*"".Func   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �<go.string.hdr."*doc.methodSet"                       4go.string."*doc.methodSet"   �4go.string."*doc.methodSet"    *doc.methodSet  �&go.string.hdr."doc"                       go.string."doc"   �go.string."doc"   doc  �2go.string.hdr."methodSet"             	          *go.string."methodSet"   �*go.string."methodSet"    methodSet  �&go.string.hdr."set"                       go.string."set"   �go.string."set"   set  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·2a1dd1e1e59d0a384c26951e316cd7e6             �&go.string.hdr."add"                       go.string."add"   �go.string."add"   add  �Tgclocals·311743cc5ea08f25d41b6a4d25949ffe 0  0                    �Tgclocals·6412d3717715814cae1af4eeac4eb5d3 0  0                   �^go.string.hdr."func(*doc.methodSet, *doc.Func)"                       Vgo.string."func(*doc.methodSet, *doc.Func)"   �Vgo.string."func(*doc.methodSet, *doc.Func)" @  @func(*doc.methodSet, *doc.Func)  �Dtype.func(*"".methodSet, *"".Func) �  �              ���f 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(*doc.methodSet, *doc.Func)"   p  Vgo.weak.type.*func(*"".methodSet, *"".Func)   �� Dtype.func(*"".methodSet, *"".Func)   �� Dtype.func(*"".methodSet, *"".Func)   �  $type.*"".methodSet   �  type.*"".Func   ��go.typelink.func(*doc.methodSet, *doc.Func)	func(*"".methodSet, *"".Func)              Dtype.func(*"".methodSet, *"".Func)   �fgo.string.hdr."func(*doc.methodSet, *ast.FuncDecl)"             #          ^go.string."func(*doc.methodSet, *ast.FuncDecl)"   �^go.string."func(*doc.methodSet, *ast.FuncDecl)" P  Hfunc(*doc.methodSet, *ast.FuncDecl)  �Ttype.func(*"".methodSet, *go/ast.FuncDecl) �  �              j�� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  fgo.string.hdr."func(*doc.methodSet, *ast.FuncDecl)"   p  fgo.weak.type.*func(*"".methodSet, *go/ast.FuncDecl)   �� Ttype.func(*"".methodSet, *go/ast.FuncDecl)   �� Ttype.func(*"".methodSet, *go/ast.FuncDecl)   �  $type.*"".methodSet   �  *type.*go/ast.FuncDecl   ��go.typelink.func(*doc.methodSet, *ast.FuncDecl)	func(*"".methodSet, *go/ast.FuncDecl)              Ttype.func(*"".methodSet, *go/ast.FuncDecl)   �>go.string.hdr."func(*doc.Func)"                       6go.string."func(*doc.Func)"   �6go.string."func(*doc.Func)"     func(*doc.Func)  �&type.func(*"".Func) �  �              מ� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."func(*doc.Func)"   p  8go.weak.type.*func(*"".Func)   �� &type.func(*"".Func)   �� &type.func(*"".Func)   �  type.*"".Func   �Tgo.typelink.func(*doc.Func)	func(*"".Func)              &type.func(*"".Func)   �Fgo.string.hdr."func(*ast.FuncDecl)"                       >go.string."func(*ast.FuncDecl)"   �>go.string."func(*ast.FuncDecl)" 0  (func(*ast.FuncDecl)  �6type.func(*go/ast.FuncDecl) �  �              � � 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."func(*ast.FuncDecl)"   p  Hgo.weak.type.*func(*go/ast.FuncDecl)   �� 6type.func(*go/ast.FuncDecl)   �� 6type.func(*go/ast.FuncDecl)   �  *type.*go/ast.FuncDecl   �lgo.typelink.func(*ast.FuncDecl)	func(*go/ast.FuncDecl)              6type.func(*go/ast.FuncDecl)   �$type.*"".methodSet  �  �              Cs�� 6                                                                                                                                                                                      &0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."*doc.methodSet"   p  6go.weak.type.**"".methodSet   �  "type."".methodSet   `� $type.*"".methodSet   �� $type.*"".methodSet   �  &go.string.hdr."add"   �  "go.importpath."".   �  &type.func(*"".Func)   �  Dtype.func(*"".methodSet, *"".Func)   �  &"".(*methodSet).add   �  &"".(*methodSet).add   �  &go.string.hdr."set"   �  "go.importpath."".   �  6type.func(*go/ast.FuncDecl)   �  Ttype.func(*"".methodSet, *go/ast.FuncDecl)   �  &"".(*methodSet).set   �  &"".(*methodSet).set   �:go.string.hdr."doc.methodSet"                       2go.string."doc.methodSet"   �2go.string."doc.methodSet"    doc.methodSet  �\go.string.hdr."func(doc.methodSet, *doc.Func)"                       Tgo.string."func(doc.methodSet, *doc.Func)"   �Tgo.string."func(doc.methodSet, *doc.Func)" @  >func(doc.methodSet, *doc.Func)  �Btype.func("".methodSet, *"".Func) �  �              �r� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(doc.methodSet, *doc.Func)"   p  Tgo.weak.type.*func("".methodSet, *"".Func)   �� Btype.func("".methodSet, *"".Func)   �� Btype.func("".methodSet, *"".Func)   �  "type."".methodSet   �  type.*"".Func   ��go.typelink.func(doc.methodSet, *doc.Func)	func("".methodSet, *"".Func)              Btype.func("".methodSet, *"".Func)   �dgo.string.hdr."func(doc.methodSet, *ast.FuncDecl)"             "          \go.string."func(doc.methodSet, *ast.FuncDecl)"   �\go.string."func(doc.methodSet, *ast.FuncDecl)" P  Ffunc(doc.methodSet, *ast.FuncDecl)  �Rtype.func("".methodSet, *go/ast.FuncDecl) �  �              w�� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  dgo.string.hdr."func(doc.methodSet, *ast.FuncDecl)"   p  dgo.weak.type.*func("".methodSet, *go/ast.FuncDecl)   �� Rtype.func("".methodSet, *go/ast.FuncDecl)   �� Rtype.func("".methodSet, *go/ast.FuncDecl)   �  "type."".methodSet   �  *type.*go/ast.FuncDecl   ��go.typelink.func(doc.methodSet, *ast.FuncDecl)	func("".methodSet, *go/ast.FuncDecl)              Rtype.func("".methodSet, *go/ast.FuncDecl)   �"type."".methodSet  �  �              C�� 5                                                                          �                                                                                                                                       00�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."doc.methodSet"   p  $type.*"".methodSet   �  type.string   �  type.*"".Func   �  >type.map.bucket[string]*"".Func   �  8type.map.hdr[string]*"".Func   `� "type."".methodSet   �  2go.string.hdr."methodSet"   �  "go.importpath."".   �� "type."".methodSet   �  &go.string.hdr."add"   �  "go.importpath."".   �  &type.func(*"".Func)   �  Btype.func("".methodSet, *"".Func)   �   "".methodSet.add   �   "".methodSet.add   �  &go.string.hdr."set"   �  "go.importpath."".   �  6type.func(*go/ast.FuncDecl)   �  Rtype.func("".methodSet, *go/ast.FuncDecl)   �   "".methodSet.set   �   "".methodSet.set   �&runtime.gcbits.d50c   � �:go.string.hdr."doc.namedType"                       2go.string."doc.namedType"   �2go.string."doc.namedType"    doc.namedType  �(go.string.hdr."name"                        go.string."name"   � go.string."name"   
name  �(go.string.hdr."decl"                        go.string."decl"   � go.string."decl"   
decl  �4go.string.hdr."isEmbedded"             
          ,go.string."isEmbedded"   �,go.string."isEmbedded"    isEmbedded  �0go.string.hdr."isStruct"                       (go.string."isStruct"   �(go.string."isStruct"    isStruct  �0go.string.hdr."embedded"                       (go.string."embedded"   �(go.string."embedded"    embedded  �*go.string.hdr."funcs"                       "go.string."funcs"   �"go.string."funcs"   funcs  �.go.string.hdr."methods"                       &go.string."methods"   �&go.string."methods"   methods  �2go.string.hdr."namedType"             	          *go.string."namedType"   �*go.string."namedType"    namedType  �"type."".namedType  �  �`       `       �7��                                                 	       	                                                                                                                                                              (                                       )                                       0                                       8                                       P                                       X                                               H0�  runtime.algarray   @  &runtime.gcbits.d50c   P  :go.string.hdr."doc.namedType"   p  $type.*"".namedType   �� "type."".namedType   �  &go.string.hdr."doc"   �  "go.importpath."".   �  type.string   �  (go.string.hdr."name"   �  "go.importpath."".   �  type.string   �  (go.string.hdr."decl"   �  "go.importpath."".   �  (type.*go/ast.GenDecl   �  4go.string.hdr."isEmbedded"   �  "go.importpath."".   �  type.bool   �  0go.string.hdr."isStruct"   �  "go.importpath."".   �  type.bool   �  0go.string.hdr."embedded"   �  "go.importpath."".   �  &type."".embeddedSet   �  ,go.string.hdr."values"   �  "go.importpath."".   �   type.[]*"".Value   �  *go.string.hdr."funcs"   �  "go.importpath."".   �  "type."".methodSet   �  .go.string.hdr."methods"   �  "go.importpath."".   �  "type."".methodSet   `� "type."".namedType   �  2go.string.hdr."namedType"   �  "go.importpath."".   �� "type."".namedType   �<go.string.hdr."*doc.namedType"                       4go.string."*doc.namedType"   �4go.string."*doc.namedType"    *doc.namedType  �$type.*"".namedType  �  �              w�� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."*doc.namedType"   p  6go.weak.type.**"".namedType   �  "type."".namedType   �bgo.string.hdr."*map.bucket[string]*doc.namedType"             !          Zgo.string."*map.bucket[string]*doc.namedType"   �Zgo.string."*map.bucket[string]*doc.namedType" P  D*map.bucket[string]*doc.namedType  �Jtype.*map.bucket[string]*"".namedType �  �              �Ny� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."*map.bucket[string]*doc.namedType"   p  \go.weak.type.**map.bucket[string]*"".namedType   �  Htype.map.bucket[string]*"".namedType   �`go.string.hdr."map.bucket[string]*doc.namedType"                        Xgo.string."map.bucket[string]*doc.namedType"   �Xgo.string."map.bucket[string]*doc.namedType" P  Bmap.bucket[string]*doc.namedType  �Htype.map.bucket[string]*"".namedType �  ��       �       �YF                                                                                                                                                                              �                                       �       0�  runtime.algarray   @  .runtime.gcbits.aaaafe03   P  `go.string.hdr."map.bucket[string]*doc.namedType"   p  Zgo.weak.type.*map.bucket[string]*"".namedType   �� Htype.map.bucket[string]*"".namedType   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  type.[8]string   �  ,go.string.hdr."values"   �  *type.[8]*"".namedType   �  0go.string.hdr."overflow"   �  Jtype.*map.bucket[string]*"".namedType   �Zgo.string.hdr."map.hdr[string]*doc.namedType"                       Rgo.string."map.hdr[string]*doc.namedType"   �Rgo.string."map.hdr[string]*doc.namedType" @  <map.hdr[string]*doc.namedType  �Btype.map.hdr[string]*"".namedType �  �0       0       $��                                                                                                                                                                              	                                                                                                                                                                                                    (       *0�  runtime.algarray   @  "runtime.gcbits.2c   P  Zgo.string.hdr."map.hdr[string]*doc.namedType"   p  Tgo.weak.type.*map.hdr[string]*"".namedType   �� Btype.map.hdr[string]*"".namedType   �  *go.string.hdr."count"   �  type.int   �  *go.string.hdr."flags"   �  type.uint8   �  "go.string.hdr."B"   �  type.uint8   �  *go.string.hdr."hash0"   �  type.uint32   �  .go.string.hdr."buckets"   �  Jtype.*map.bucket[string]*"".namedType   �  4go.string.hdr."oldbuckets"   �  Jtype.*map.bucket[string]*"".namedType   �  2go.string.hdr."nevacuate"   �  type.uintptr   �  0go.string.hdr."overflow"   �  &type.unsafe.Pointer   �Rgo.string.hdr."map[string]*doc.namedType"                       Jgo.string."map[string]*doc.namedType"   �Jgo.string."map[string]*doc.namedType" @  4map[string]*doc.namedType  �:type.map[string]*"".namedType �  �              ��� 5                                                                          � 0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."map[string]*doc.namedType"   p  Lgo.weak.type.*map[string]*"".namedType   �  type.string   �  $type.*"".namedType   �  Htype.map.bucket[string]*"".namedType   �  Btype.map.hdr[string]*"".namedType   �|go.typelink.map[string]*doc.namedType	map[string]*"".namedType              :type.map[string]*"".namedType   �Hgo.string.hdr."[]*ast.InterfaceType"                       @go.string."[]*ast.InterfaceType"   �@go.string."[]*ast.InterfaceType" 0  *[]*ast.InterfaceType  �8type.[]*go/ast.InterfaceType �  �              �b�-                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."[]*ast.InterfaceType"   p  Jgo.weak.type.*[]*go/ast.InterfaceType   �  4type.*go/ast.InterfaceType   �pgo.typelink.[]*ast.InterfaceType	[]*go/ast.InterfaceType              8type.[]*go/ast.InterfaceType   �6go.string.hdr."*doc.reader"                       .go.string."*doc.reader"   �.go.string."*doc.reader"    *doc.reader  �Bgo.string.hdr."func(*doc.reader)"                       :go.string."func(*doc.reader)"   �:go.string."func(*doc.reader)" 0  $func(*doc.reader)  �*type.func(*"".reader) �  �              �Ik 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."func(*doc.reader)"   p  <go.weak.type.*func(*"".reader)   �� *type.func(*"".reader)   �� *type.func(*"".reader)   �  type.*"".reader   �\go.typelink.func(*doc.reader)	func(*"".reader)              *type.func(*"".reader)   ��go.string.hdr."func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"             T          �go.string."func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"   ��go.string."func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)" �  �func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)  ��type.func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet) �  �              �0$d 3                                                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"   p  �go.weak.type.*func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �� �type.func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �� �type.func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �  type.*"".reader   �  "type."".methodSet   �  $type.*"".namedType   �  type.string   �  type.bool   �  type.int   �  &type."".embeddedSet   ��go.typelink.func(*doc.reader, doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)	func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)              �type.func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �Xgo.string.hdr."func(*doc.reader, *ast.File)"                       Pgo.string."func(*doc.reader, *ast.File)"   �Pgo.string."func(*doc.reader, *ast.File)" @  :func(*doc.reader, *ast.File)  �Ftype.func(*"".reader, *go/ast.File) �  �              �+( 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."func(*doc.reader, *ast.File)"   p  Xgo.weak.type.*func(*"".reader, *go/ast.File)   �� Ftype.func(*"".reader, *go/ast.File)   �� Ftype.func(*"".reader, *go/ast.File)   �  type.*"".reader   �  "type.*go/ast.File   ��go.typelink.func(*doc.reader, *ast.File)	func(*"".reader, *go/ast.File)              Ftype.func(*"".reader, *go/ast.File)   �`go.string.hdr."func(*doc.reader, ast.Decl) bool"                        Xgo.string."func(*doc.reader, ast.Decl) bool"   �Xgo.string."func(*doc.reader, ast.Decl) bool" P  Bfunc(*doc.reader, ast.Decl) bool  �Ntype.func(*"".reader, go/ast.Decl) bool �  �              "�+ 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(*doc.reader, ast.Decl) bool"   p  `go.weak.type.*func(*"".reader, go/ast.Decl) bool   �� Ntype.func(*"".reader, go/ast.Decl) bool   �� Ntype.func(*"".reader, go/ast.Decl) bool   �  type.*"".reader   �   type.go/ast.Decl   �  type.bool   ��go.typelink.func(*doc.reader, ast.Decl) bool	func(*"".reader, go/ast.Decl) bool              Ntype.func(*"".reader, go/ast.Decl) bool   ��go.string.hdr."func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"             J          �go.string."func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"   ��go.string."func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool" �  �func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool  ��type.func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool �  �              ��$� 3                                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"   p  �go.weak.type.*func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �� �type.func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �� �type.func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �  type.*"".reader   �  $type.*"".namedType   �  ,type.*go/ast.FieldList   �  4type.*go/ast.InterfaceType   �  type.bool   ��go.typelink.func(*doc.reader, *doc.namedType, *ast.FieldList, *ast.InterfaceType) bool	func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool              �type.func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �bgo.string.hdr."func(*doc.reader, *ast.FieldList)"             !          Zgo.string."func(*doc.reader, *ast.FieldList)"   �Zgo.string."func(*doc.reader, *ast.FieldList)" P  Dfunc(*doc.reader, *ast.FieldList)  �Ptype.func(*"".reader, *go/ast.FieldList) �  �              (��� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*doc.reader, *ast.FieldList)"   p  bgo.weak.type.*func(*"".reader, *go/ast.FieldList)   �� Ptype.func(*"".reader, *go/ast.FieldList)   �� Ptype.func(*"".reader, *go/ast.FieldList)   �  type.*"".reader   �  ,type.*go/ast.FieldList   ��go.typelink.func(*doc.reader, *ast.FieldList)	func(*"".reader, *go/ast.FieldList)              Ptype.func(*"".reader, *go/ast.FieldList)   �zgo.string.hdr."func(*doc.reader, ast.Spec, token.Token) bool"             -          rgo.string."func(*doc.reader, ast.Spec, token.Token) bool"   �rgo.string."func(*doc.reader, ast.Spec, token.Token) bool" `  \func(*doc.reader, ast.Spec, token.Token) bool  �ntype.func(*"".reader, go/ast.Spec, go/token.Token) bool �  �              B�* 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  zgo.string.hdr."func(*doc.reader, ast.Spec, token.Token) bool"   p  �go.weak.type.*func(*"".reader, go/ast.Spec, go/token.Token) bool   �� ntype.func(*"".reader, go/ast.Spec, go/token.Token) bool   �� ntype.func(*"".reader, go/ast.Spec, go/token.Token) bool   �  type.*"".reader   �   type.go/ast.Spec   �  &type.go/token.Token   �  type.bool   ��go.typelink.func(*doc.reader, ast.Spec, token.Token) bool	func(*"".reader, go/ast.Spec, go/token.Token) bool              ntype.func(*"".reader, go/ast.Spec, go/token.Token) bool   �4go.string.hdr."[]ast.Spec"             
          ,go.string."[]ast.Spec"   �,go.string."[]ast.Spec"    []ast.Spec  �$type.[]go/ast.Spec �  �              0�4                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."[]ast.Spec"   p  6go.weak.type.*[]go/ast.Spec   �   type.go/ast.Spec   �Hgo.typelink.[]ast.Spec	[]go/ast.Spec              $type.[]go/ast.Spec   ��go.string.hdr."func(*doc.reader, []ast.Spec, token.Token) []ast.Spec"             5          �go.string."func(*doc.reader, []ast.Spec, token.Token) []ast.Spec"   ��go.string."func(*doc.reader, []ast.Spec, token.Token) []ast.Spec" p  lfunc(*doc.reader, []ast.Spec, token.Token) []ast.Spec  ��type.func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec �  �              /=� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*doc.reader, []ast.Spec, token.Token) []ast.Spec"   p  �go.weak.type.*func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec   �� �type.func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec   �� �type.func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec   �  type.*"".reader   �  $type.[]go/ast.Spec   �  &type.go/token.Token   �  $type.[]go/ast.Spec   ��go.typelink.func(*doc.reader, []ast.Spec, token.Token) []ast.Spec	func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec              �type.func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec   �vgo.string.hdr."func(*doc.reader, *doc.namedType, ast.Expr)"             +          ngo.string."func(*doc.reader, *doc.namedType, ast.Expr)"   �ngo.string."func(*doc.reader, *doc.namedType, ast.Expr)" `  Xfunc(*doc.reader, *doc.namedType, ast.Expr)  �btype.func(*"".reader, *"".namedType, go/ast.Expr) �  �              �e�� 3                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  vgo.string.hdr."func(*doc.reader, *doc.namedType, ast.Expr)"   p  tgo.weak.type.*func(*"".reader, *"".namedType, go/ast.Expr)   �� btype.func(*"".reader, *"".namedType, go/ast.Expr)   �� btype.func(*"".reader, *"".namedType, go/ast.Expr)   �  type.*"".reader   �  $type.*"".namedType   �   type.go/ast.Expr   ��go.typelink.func(*doc.reader, *doc.namedType, ast.Expr)	func(*"".reader, *"".namedType, go/ast.Expr)              btype.func(*"".reader, *"".namedType, go/ast.Expr)   �\go.string.hdr."func(*doc.reader, string) bool"                       Tgo.string."func(*doc.reader, string) bool"   �Tgo.string."func(*doc.reader, string) bool" @  >func(*doc.reader, string) bool  �Dtype.func(*"".reader, string) bool �  �              ��� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(*doc.reader, string) bool"   p  Vgo.weak.type.*func(*"".reader, string) bool   �� Dtype.func(*"".reader, string) bool   �� Dtype.func(*"".reader, string) bool   �  type.*"".reader   �  type.string   �  type.bool   ��go.typelink.func(*doc.reader, string) bool	func(*"".reader, string) bool              Dtype.func(*"".reader, string) bool   �pgo.string.hdr."func(*doc.reader, string) *doc.namedType"             (          hgo.string."func(*doc.reader, string) *doc.namedType"   �hgo.string."func(*doc.reader, string) *doc.namedType" `  Rfunc(*doc.reader, string) *doc.namedType  �Vtype.func(*"".reader, string) *"".namedType �  �              [52 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  pgo.string.hdr."func(*doc.reader, string) *doc.namedType"   p  hgo.weak.type.*func(*"".reader, string) *"".namedType   �� Vtype.func(*"".reader, string) *"".namedType   �� Vtype.func(*"".reader, string) *"".namedType   �  type.*"".reader   �  type.string   �  $type.*"".namedType   ��go.typelink.func(*doc.reader, string) *doc.namedType	func(*"".reader, string) *"".namedType              Vtype.func(*"".reader, string) *"".namedType   �hgo.string.hdr."func(*doc.reader, *ast.CommentGroup)"             $          `go.string."func(*doc.reader, *ast.CommentGroup)"   �`go.string."func(*doc.reader, *ast.CommentGroup)" P  Jfunc(*doc.reader, *ast.CommentGroup)  �Vtype.func(*"".reader, *go/ast.CommentGroup) �  �              �vl 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  hgo.string.hdr."func(*doc.reader, *ast.CommentGroup)"   p  hgo.weak.type.*func(*"".reader, *go/ast.CommentGroup)   �� Vtype.func(*"".reader, *go/ast.CommentGroup)   �� Vtype.func(*"".reader, *go/ast.CommentGroup)   �  type.*"".reader   �  2type.*go/ast.CommentGroup   ��go.typelink.func(*doc.reader, *ast.CommentGroup)	func(*"".reader, *go/ast.CommentGroup)              Vtype.func(*"".reader, *go/ast.CommentGroup)   �`go.string.hdr."func(*doc.reader, *ast.FuncDecl)"                        Xgo.string."func(*doc.reader, *ast.FuncDecl)"   �Xgo.string."func(*doc.reader, *ast.FuncDecl)" P  Bfunc(*doc.reader, *ast.FuncDecl)  �Ntype.func(*"".reader, *go/ast.FuncDecl) �  �              �A�� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(*doc.reader, *ast.FuncDecl)"   p  `go.weak.type.*func(*"".reader, *go/ast.FuncDecl)   �� Ntype.func(*"".reader, *go/ast.FuncDecl)   �� Ntype.func(*"".reader, *go/ast.FuncDecl)   �  type.*"".reader   �  *type.*go/ast.FuncDecl   ��go.typelink.func(*doc.reader, *ast.FuncDecl)	func(*"".reader, *go/ast.FuncDecl)              Ntype.func(*"".reader, *go/ast.FuncDecl)   �<go.string.hdr."[]*ast.Comment"                       4go.string."[]*ast.Comment"   �4go.string."[]*ast.Comment"    []*ast.Comment  �,type.[]*go/ast.Comment �  �              5~�                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."[]*ast.Comment"   p  >go.weak.type.*[]*go/ast.Comment   �  (type.*go/ast.Comment   �Xgo.typelink.[]*ast.Comment	[]*go/ast.Comment              ,type.[]*go/ast.Comment   �bgo.string.hdr."func(*doc.reader, []*ast.Comment)"             !          Zgo.string."func(*doc.reader, []*ast.Comment)"   �Zgo.string."func(*doc.reader, []*ast.Comment)" P  Dfunc(*doc.reader, []*ast.Comment)  �Ptype.func(*"".reader, []*go/ast.Comment) �  �              E@5i 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*doc.reader, []*ast.Comment)"   p  bgo.weak.type.*func(*"".reader, []*go/ast.Comment)   �� Ptype.func(*"".reader, []*go/ast.Comment)   �� Ptype.func(*"".reader, []*go/ast.Comment)   �  type.*"".reader   �  ,type.[]*go/ast.Comment   ��go.typelink.func(*doc.reader, []*ast.Comment)	func(*"".reader, []*go/ast.Comment)              Ptype.func(*"".reader, []*go/ast.Comment)   �Fgo.string.hdr."[]*ast.CommentGroup"                       >go.string."[]*ast.CommentGroup"   �>go.string."[]*ast.CommentGroup" 0  ([]*ast.CommentGroup  �6type.[]*go/ast.CommentGroup �  �              �b�i                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."[]*ast.CommentGroup"   p  Hgo.weak.type.*[]*go/ast.CommentGroup   �  2type.*go/ast.CommentGroup   �lgo.typelink.[]*ast.CommentGroup	[]*go/ast.CommentGroup              6type.[]*go/ast.CommentGroup   �lgo.string.hdr."func(*doc.reader, []*ast.CommentGroup)"             &          dgo.string."func(*doc.reader, []*ast.CommentGroup)"   �dgo.string."func(*doc.reader, []*ast.CommentGroup)" P  Nfunc(*doc.reader, []*ast.CommentGroup)  �Ztype.func(*"".reader, []*go/ast.CommentGroup) �  �              ��� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(*doc.reader, []*ast.CommentGroup)"   p  lgo.weak.type.*func(*"".reader, []*go/ast.CommentGroup)   �� Ztype.func(*"".reader, []*go/ast.CommentGroup)   �� Ztype.func(*"".reader, []*go/ast.CommentGroup)   �  type.*"".reader   �  6type.[]*go/ast.CommentGroup   ��go.typelink.func(*doc.reader, []*ast.CommentGroup)	func(*"".reader, []*go/ast.CommentGroup)              Ztype.func(*"".reader, []*go/ast.CommentGroup)   �rgo.string.hdr."func(*doc.reader, *ast.Package, doc.Mode)"             )          jgo.string."func(*doc.reader, *ast.Package, doc.Mode)"   �jgo.string."func(*doc.reader, *ast.Package, doc.Mode)" `  Tfunc(*doc.reader, *ast.Package, doc.Mode)  �^type.func(*"".reader, *go/ast.Package, "".Mode) �  �              <Pt� 3                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  rgo.string.hdr."func(*doc.reader, *ast.Package, doc.Mode)"   p  pgo.weak.type.*func(*"".reader, *go/ast.Package, "".Mode)   �� ^type.func(*"".reader, *go/ast.Package, "".Mode)   �� ^type.func(*"".reader, *go/ast.Package, "".Mode)   �  type.*"".reader   �  (type.*go/ast.Package   �  type."".Mode   ��go.typelink.func(*doc.reader, *ast.Package, doc.Mode)	func(*"".reader, *go/ast.Package, "".Mode)              ^type.func(*"".reader, *go/ast.Package, "".Mode)   �|go.string.hdr."func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)"             .          tgo.string."func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)"   �tgo.string."func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)" `  ^func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)  �ptype.func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec) �  �              �2 3                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  |go.string.hdr."func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)"   p  �go.weak.type.*func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)   �� ptype.func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)   �� ptype.func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)   �  type.*"".reader   �  (type.*go/ast.GenDecl   �  *type.*go/ast.TypeSpec   ��go.typelink.func(*doc.reader, *ast.GenDecl, *ast.TypeSpec)	func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)              ptype.func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)   �^go.string.hdr."func(*doc.reader, *ast.GenDecl)"                       Vgo.string."func(*doc.reader, *ast.GenDecl)"   �Vgo.string."func(*doc.reader, *ast.GenDecl)" @  @func(*doc.reader, *ast.GenDecl)  �Ltype.func(*"".reader, *go/ast.GenDecl) �  �              �&V 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  ^go.string.hdr."func(*doc.reader, *ast.GenDecl)"   p  ^go.weak.type.*func(*"".reader, *go/ast.GenDecl)   �� Ltype.func(*"".reader, *go/ast.GenDecl)   �� Ltype.func(*"".reader, *go/ast.GenDecl)   �  type.*"".reader   �  (type.*go/ast.GenDecl   ��go.typelink.func(*doc.reader, *ast.GenDecl)	func(*"".reader, *go/ast.GenDecl)              Ltype.func(*"".reader, *go/ast.GenDecl)   ��go.string.hdr."func(*doc.reader, *doc.namedType, ast.Expr) string"             2          |go.string."func(*doc.reader, *doc.namedType, ast.Expr) string"   �|go.string."func(*doc.reader, *doc.namedType, ast.Expr) string" p  ffunc(*doc.reader, *doc.namedType, ast.Expr) string  �ptype.func(*"".reader, *"".namedType, go/ast.Expr) string �  �              �
�{ 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*doc.reader, *doc.namedType, ast.Expr) string"   p  �go.weak.type.*func(*"".reader, *"".namedType, go/ast.Expr) string   �� ptype.func(*"".reader, *"".namedType, go/ast.Expr) string   �� ptype.func(*"".reader, *"".namedType, go/ast.Expr) string   �  type.*"".reader   �  $type.*"".namedType   �   type.go/ast.Expr   �  type.string   ��go.typelink.func(*doc.reader, *doc.namedType, ast.Expr) string	func(*"".reader, *"".namedType, go/ast.Expr) string              ptype.func(*"".reader, *"".namedType, go/ast.Expr) string   �jgo.string.hdr."func(*doc.reader, *ast.InterfaceType)"             %          bgo.string."func(*doc.reader, *ast.InterfaceType)"   �bgo.string."func(*doc.reader, *ast.InterfaceType)" P  Lfunc(*doc.reader, *ast.InterfaceType)  �Xtype.func(*"".reader, *go/ast.InterfaceType) �  �              �}� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(*doc.reader, *ast.InterfaceType)"   p  jgo.weak.type.*func(*"".reader, *go/ast.InterfaceType)   �� Xtype.func(*"".reader, *go/ast.InterfaceType)   �� Xtype.func(*"".reader, *go/ast.InterfaceType)   �  type.*"".reader   �  4type.*go/ast.InterfaceType   ��go.typelink.func(*doc.reader, *ast.InterfaceType)	func(*"".reader, *go/ast.InterfaceType)              Xtype.func(*"".reader, *go/ast.InterfaceType)   �8go.string.hdr."cleanupTypes"                       0go.string."cleanupTypes"   �0go.string."cleanupTypes"    cleanupTypes  �Lgo.string.hdr."collectEmbeddedMethods"                       Dgo.string."collectEmbeddedMethods"   �Dgo.string."collectEmbeddedMethods" 0  .collectEmbeddedMethods  ��go.string.hdr."func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"             G          �go.string."func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"   ��go.string."func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)" �  �func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)  ��type.func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet) �  �              ʦ�X 3                                                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)"   p  �go.weak.type.*func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �� �type.func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �� �type.func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �  "type."".methodSet   �  $type.*"".namedType   �  type.string   �  type.bool   �  type.int   �  &type."".embeddedSet   ��go.typelink.func(doc.methodSet, *doc.namedType, string, bool, int, doc.embeddedSet)	func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)              �type.func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �Bgo.string.hdr."computeMethodSets"                       :go.string."computeMethodSets"   �:go.string."computeMethodSets" 0  $computeMethodSets  �6go.string.hdr."fileExports"                       .go.string."fileExports"   �.go.string."fileExports"    fileExports  �>go.string.hdr."func(*ast.File)"                       6go.string."func(*ast.File)"   �6go.string."func(*ast.File)"     func(*ast.File)  �.type.func(*go/ast.File) �  �              �~K 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  >go.string.hdr."func(*ast.File)"   p  @go.weak.type.*func(*go/ast.File)   �� .type.func(*go/ast.File)   �� .type.func(*go/ast.File)   �  "type.*go/ast.File   �\go.typelink.func(*ast.File)	func(*go/ast.File)              .type.func(*go/ast.File)   �4go.string.hdr."filterDecl"             
          ,go.string."filterDecl"   �,go.string."filterDecl"    filterDecl  �Fgo.string.hdr."func(ast.Decl) bool"                       >go.string."func(ast.Decl) bool"   �>go.string."func(ast.Decl) bool" 0  (func(ast.Decl) bool  �6type.func(go/ast.Decl) bool �  �              �j�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."func(ast.Decl) bool"   p  Hgo.weak.type.*func(go/ast.Decl) bool   �� 6type.func(go/ast.Decl) bool   �� 6type.func(go/ast.Decl) bool   �   type.go/ast.Decl   �  type.bool   �lgo.typelink.func(ast.Decl) bool	func(go/ast.Decl) bool              6type.func(go/ast.Decl) bool   �>go.string.hdr."filterFieldList"                       6go.string."filterFieldList"   �6go.string."filterFieldList"     filterFieldList  ��go.string.hdr."func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"             =          �go.string."func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"   ��go.string."func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool" �  |func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool  ��type.func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool �  �              �� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  �go.string.hdr."func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool"   p  �go.weak.type.*func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �� �type.func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �� �type.func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �  $type.*"".namedType   �  ,type.*go/ast.FieldList   �  4type.*go/ast.InterfaceType   �  type.bool   ��go.typelink.func(*doc.namedType, *ast.FieldList, *ast.InterfaceType) bool	func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool              �type.func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �>go.string.hdr."filterParamList"                       6go.string."filterParamList"   �6go.string."filterParamList"     filterParamList  �Hgo.string.hdr."func(*ast.FieldList)"                       @go.string."func(*ast.FieldList)"   �@go.string."func(*ast.FieldList)" 0  *func(*ast.FieldList)  �8type.func(*go/ast.FieldList) �  �              x/� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."func(*ast.FieldList)"   p  Jgo.weak.type.*func(*go/ast.FieldList)   �� 8type.func(*go/ast.FieldList)   �� 8type.func(*go/ast.FieldList)   �  ,type.*go/ast.FieldList   �pgo.typelink.func(*ast.FieldList)	func(*go/ast.FieldList)              8type.func(*go/ast.FieldList)   �4go.string.hdr."filterSpec"             
          ,go.string."filterSpec"   �,go.string."filterSpec"    filterSpec  �`go.string.hdr."func(ast.Spec, token.Token) bool"                        Xgo.string."func(ast.Spec, token.Token) bool"   �Xgo.string."func(ast.Spec, token.Token) bool" P  Bfunc(ast.Spec, token.Token) bool  �Vtype.func(go/ast.Spec, go/token.Token) bool �  �              �G�� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  `go.string.hdr."func(ast.Spec, token.Token) bool"   p  hgo.weak.type.*func(go/ast.Spec, go/token.Token) bool   �� Vtype.func(go/ast.Spec, go/token.Token) bool   �� Vtype.func(go/ast.Spec, go/token.Token) bool   �   type.go/ast.Spec   �  &type.go/token.Token   �  type.bool   ��go.typelink.func(ast.Spec, token.Token) bool	func(go/ast.Spec, go/token.Token) bool              Vtype.func(go/ast.Spec, go/token.Token) bool   �<go.string.hdr."filterSpecList"                       4go.string."filterSpecList"   �4go.string."filterSpecList"    filterSpecList  �pgo.string.hdr."func([]ast.Spec, token.Token) []ast.Spec"             (          hgo.string."func([]ast.Spec, token.Token) []ast.Spec"   �hgo.string."func([]ast.Spec, token.Token) []ast.Spec" `  Rfunc([]ast.Spec, token.Token) []ast.Spec  �ltype.func([]go/ast.Spec, go/token.Token) []go/ast.Spec �  �              �\
 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  pgo.string.hdr."func([]ast.Spec, token.Token) []ast.Spec"   p  ~go.weak.type.*func([]go/ast.Spec, go/token.Token) []go/ast.Spec   �� ltype.func([]go/ast.Spec, go/token.Token) []go/ast.Spec   �� ltype.func([]go/ast.Spec, go/token.Token) []go/ast.Spec   �  $type.[]go/ast.Spec   �  &type.go/token.Token   �  $type.[]go/ast.Spec   ��go.typelink.func([]ast.Spec, token.Token) []ast.Spec	func([]go/ast.Spec, go/token.Token) []go/ast.Spec              ltype.func([]go/ast.Spec, go/token.Token) []go/ast.Spec   �4go.string.hdr."filterType"             
          ,go.string."filterType"   �,go.string."filterType"    filterType  �\go.string.hdr."func(*doc.namedType, ast.Expr)"                       Tgo.string."func(*doc.namedType, ast.Expr)"   �Tgo.string."func(*doc.namedType, ast.Expr)" @  >func(*doc.namedType, ast.Expr)  �Jtype.func(*"".namedType, go/ast.Expr) �  �              գ�� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  \go.string.hdr."func(*doc.namedType, ast.Expr)"   p  \go.weak.type.*func(*"".namedType, go/ast.Expr)   �� Jtype.func(*"".namedType, go/ast.Expr)   �� Jtype.func(*"".namedType, go/ast.Expr)   �  $type.*"".namedType   �   type.go/ast.Expr   ��go.typelink.func(*doc.namedType, ast.Expr)	func(*"".namedType, go/ast.Expr)              Jtype.func(*"".namedType, go/ast.Expr)   �2go.string.hdr."isVisible"             	          *go.string."isVisible"   �*go.string."isVisible"    isVisible  �Bgo.string.hdr."func(string) bool"                       :go.string."func(string) bool"   �:go.string."func(string) bool" 0  $func(string) bool  �,type.func(string) bool �  �              *�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."func(string) bool"   p  >go.weak.type.*func(string) bool   �� ,type.func(string) bool   �� ,type.func(string) bool   �  type.string   �  type.bool   �^go.typelink.func(string) bool	func(string) bool              ,type.func(string) bool   �4go.string.hdr."lookupType"             
          ,go.string."lookupType"   �,go.string."lookupType"    lookupType  �Vgo.string.hdr."func(string) *doc.namedType"                       Ngo.string."func(string) *doc.namedType"   �Ngo.string."func(string) *doc.namedType" @  8func(string) *doc.namedType  �>type.func(string) *"".namedType �  �              M
 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Vgo.string.hdr."func(string) *doc.namedType"   p  Pgo.weak.type.*func(string) *"".namedType   �� >type.func(string) *"".namedType   �� >type.func(string) *"".namedType   �  type.string   �  $type.*"".namedType   ��go.typelink.func(string) *doc.namedType	func(string) *"".namedType              >type.func(string) *"".namedType   �.go.string.hdr."readDoc"                       &go.string."readDoc"   �&go.string."readDoc"   readDoc  �Ngo.string.hdr."func(*ast.CommentGroup)"                       Fgo.string."func(*ast.CommentGroup)"   �Fgo.string."func(*ast.CommentGroup)" 0  0func(*ast.CommentGroup)  �>type.func(*go/ast.CommentGroup) �  �              F� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Ngo.string.hdr."func(*ast.CommentGroup)"   p  Pgo.weak.type.*func(*go/ast.CommentGroup)   �� >type.func(*go/ast.CommentGroup)   �� >type.func(*go/ast.CommentGroup)   �  2type.*go/ast.CommentGroup   �|go.typelink.func(*ast.CommentGroup)	func(*go/ast.CommentGroup)              >type.func(*go/ast.CommentGroup)   �0go.string.hdr."readFile"                       (go.string."readFile"   �(go.string."readFile"    readFile  �0go.string.hdr."readFunc"                       (go.string."readFunc"   �(go.string."readFunc"    readFunc  �0go.string.hdr."readNote"                       (go.string."readNote"   �(go.string."readNote"    readNote  �Hgo.string.hdr."func([]*ast.Comment)"                       @go.string."func([]*ast.Comment)"   �@go.string."func([]*ast.Comment)" 0  *func([]*ast.Comment)  �8type.func([]*go/ast.Comment) �  �              !� y 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Hgo.string.hdr."func([]*ast.Comment)"   p  Jgo.weak.type.*func([]*go/ast.Comment)   �� 8type.func([]*go/ast.Comment)   �� 8type.func([]*go/ast.Comment)   �  ,type.[]*go/ast.Comment   �pgo.typelink.func([]*ast.Comment)	func([]*go/ast.Comment)              8type.func([]*go/ast.Comment)   �2go.string.hdr."readNotes"             	          *go.string."readNotes"   �*go.string."readNotes"    readNotes  �Rgo.string.hdr."func([]*ast.CommentGroup)"                       Jgo.string."func([]*ast.CommentGroup)"   �Jgo.string."func([]*ast.CommentGroup)" @  4func([]*ast.CommentGroup)  �Btype.func([]*go/ast.CommentGroup) �  �              ��� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Rgo.string.hdr."func([]*ast.CommentGroup)"   p  Tgo.weak.type.*func([]*go/ast.CommentGroup)   �� Btype.func([]*go/ast.CommentGroup)   �� Btype.func([]*go/ast.CommentGroup)   �  6type.[]*go/ast.CommentGroup   ��go.typelink.func([]*ast.CommentGroup)	func([]*go/ast.CommentGroup)              Btype.func([]*go/ast.CommentGroup)   �6go.string.hdr."readPackage"                       .go.string."readPackage"   �.go.string."readPackage"    readPackage  �Xgo.string.hdr."func(*ast.Package, doc.Mode)"                       Pgo.string."func(*ast.Package, doc.Mode)"   �Pgo.string."func(*ast.Package, doc.Mode)" @  :func(*ast.Package, doc.Mode)  �Ftype.func(*go/ast.Package, "".Mode) �  �              F�m= 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."func(*ast.Package, doc.Mode)"   p  Xgo.weak.type.*func(*go/ast.Package, "".Mode)   �� Ftype.func(*go/ast.Package, "".Mode)   �� Ftype.func(*go/ast.Package, "".Mode)   �  (type.*go/ast.Package   �  type."".Mode   ��go.typelink.func(*ast.Package, doc.Mode)	func(*go/ast.Package, "".Mode)              Ftype.func(*go/ast.Package, "".Mode)   �0go.string.hdr."readType"                       (go.string."readType"   �(go.string."readType"    readType  �bgo.string.hdr."func(*ast.GenDecl, *ast.TypeSpec)"             !          Zgo.string."func(*ast.GenDecl, *ast.TypeSpec)"   �Zgo.string."func(*ast.GenDecl, *ast.TypeSpec)" P  Dfunc(*ast.GenDecl, *ast.TypeSpec)  �Xtype.func(*go/ast.GenDecl, *go/ast.TypeSpec) �  �              ŗ�� 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(*ast.GenDecl, *ast.TypeSpec)"   p  jgo.weak.type.*func(*go/ast.GenDecl, *go/ast.TypeSpec)   �� Xtype.func(*go/ast.GenDecl, *go/ast.TypeSpec)   �� Xtype.func(*go/ast.GenDecl, *go/ast.TypeSpec)   �  (type.*go/ast.GenDecl   �  *type.*go/ast.TypeSpec   ��go.typelink.func(*ast.GenDecl, *ast.TypeSpec)	func(*go/ast.GenDecl, *go/ast.TypeSpec)              Xtype.func(*go/ast.GenDecl, *go/ast.TypeSpec)   �2go.string.hdr."readValue"             	          *go.string."readValue"   �*go.string."readValue"    readValue  �Dgo.string.hdr."func(*ast.GenDecl)"                       <go.string."func(*ast.GenDecl)"   �<go.string."func(*ast.GenDecl)" 0  &func(*ast.GenDecl)  �4type.func(*go/ast.GenDecl) �  �              �^�� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."func(*ast.GenDecl)"   p  Fgo.weak.type.*func(*go/ast.GenDecl)   �� 4type.func(*go/ast.GenDecl)   �� 4type.func(*go/ast.GenDecl)   �  (type.*go/ast.GenDecl   �hgo.typelink.func(*ast.GenDecl)	func(*go/ast.GenDecl)              4type.func(*go/ast.GenDecl)   �Hgo.string.hdr."recordAnonymousField"                       @go.string."recordAnonymousField"   �@go.string."recordAnonymousField" 0  *recordAnonymousField  �jgo.string.hdr."func(*doc.namedType, ast.Expr) string"             %          bgo.string."func(*doc.namedType, ast.Expr) string"   �bgo.string."func(*doc.namedType, ast.Expr) string" P  Lfunc(*doc.namedType, ast.Expr) string  �Xtype.func(*"".namedType, go/ast.Expr) string �  �              �&� 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  jgo.string.hdr."func(*doc.namedType, ast.Expr) string"   p  jgo.weak.type.*func(*"".namedType, go/ast.Expr) string   �� Xtype.func(*"".namedType, go/ast.Expr) string   �� Xtype.func(*"".namedType, go/ast.Expr) string   �  $type.*"".namedType   �   type.go/ast.Expr   �  type.string   ��go.typelink.func(*doc.namedType, ast.Expr) string	func(*"".namedType, go/ast.Expr) string              Xtype.func(*"".namedType, go/ast.Expr) string   �0go.string.hdr."remember"                       (go.string."remember"   �(go.string."remember"    remember  �Pgo.string.hdr."func(*ast.InterfaceType)"                       Hgo.string."func(*ast.InterfaceType)"   �Hgo.string."func(*ast.InterfaceType)" @  2func(*ast.InterfaceType)  �@type.func(*go/ast.InterfaceType) �  �              x9�� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  Pgo.string.hdr."func(*ast.InterfaceType)"   p  Rgo.weak.type.*func(*go/ast.InterfaceType)   �� @type.func(*go/ast.InterfaceType)   �� @type.func(*go/ast.InterfaceType)   �  4type.*go/ast.InterfaceType   ��go.typelink.func(*ast.InterfaceType)	func(*go/ast.InterfaceType)              @type.func(*go/ast.InterfaceType)   �type.*"".reader  �  �              �}`� 6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."*doc.reader"   p  0go.weak.type.**"".reader   �  type."".reader   `� type.*"".reader   �� type.*"".reader   �  8go.string.hdr."cleanupTypes"   �  "go.importpath."".   �  type.func()   �  *type.func(*"".reader)   �  2"".(*reader).cleanupTypes   �  2"".(*reader).cleanupTypes   �  Lgo.string.hdr."collectEmbeddedMethods"   �  "go.importpath."".   �  �type.func("".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �  �type.func(*"".reader, "".methodSet, *"".namedType, string, bool, int, "".embeddedSet)   �  F"".(*reader).collectEmbeddedMethods   �  F"".(*reader).collectEmbeddedMethods   �  Bgo.string.hdr."computeMethodSets"   �  "go.importpath."".   �  type.func()   �  *type.func(*"".reader)   �  <"".(*reader).computeMethodSets   �  <"".(*reader).computeMethodSets   �  6go.string.hdr."fileExports"   �  "go.importpath."".   �  .type.func(*go/ast.File)   �  Ftype.func(*"".reader, *go/ast.File)   �  0"".(*reader).fileExports   �  0"".(*reader).fileExports   �  4go.string.hdr."filterDecl"   �  "go.importpath."".   �  6type.func(go/ast.Decl) bool   �  Ntype.func(*"".reader, go/ast.Decl) bool   �  ."".(*reader).filterDecl   �  ."".(*reader).filterDecl   �  >go.string.hdr."filterFieldList"   �  "go.importpath."".   �  �type.func(*"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �  �type.func(*"".reader, *"".namedType, *go/ast.FieldList, *go/ast.InterfaceType) bool   �  8"".(*reader).filterFieldList   �  8"".(*reader).filterFieldList   �  >go.string.hdr."filterParamList"   �  "go.importpath."".   �  8type.func(*go/ast.FieldList)   �  Ptype.func(*"".reader, *go/ast.FieldList)   �  8"".(*reader).filterParamList   �  8"".(*reader).filterParamList   �  4go.string.hdr."filterSpec"   �  "go.importpath."".   �  Vtype.func(go/ast.Spec, go/token.Token) bool   �  ntype.func(*"".reader, go/ast.Spec, go/token.Token) bool   �  ."".(*reader).filterSpec   �  ."".(*reader).filterSpec   �  <go.string.hdr."filterSpecList"   �  "go.importpath."".   �  ltype.func([]go/ast.Spec, go/token.Token) []go/ast.Spec   �  �type.func(*"".reader, []go/ast.Spec, go/token.Token) []go/ast.Spec   �  6"".(*reader).filterSpecList   �  6"".(*reader).filterSpecList   �  4go.string.hdr."filterType"   �  "go.importpath."".   �  Jtype.func(*"".namedType, go/ast.Expr)   �  btype.func(*"".reader, *"".namedType, go/ast.Expr)   �	  ."".(*reader).filterType   �	  ."".(*reader).filterType   �	  2go.string.hdr."isVisible"   �	  "go.importpath."".   �	  ,type.func(string) bool   �	  Dtype.func(*"".reader, string) bool   �	  ,"".(*reader).isVisible   �	  ,"".(*reader).isVisible   �
  4go.string.hdr."lookupType"   �
  "go.importpath."".   �
  >type.func(string) *"".namedType   �
  Vtype.func(*"".reader, string) *"".namedType   �
  ."".(*reader).lookupType   �
  ."".(*reader).lookupType   �
  .go.string.hdr."readDoc"   �
  "go.importpath."".   �  >type.func(*go/ast.CommentGroup)   �  Vtype.func(*"".reader, *go/ast.CommentGroup)   �  ("".(*reader).readDoc   �  ("".(*reader).readDoc   �  0go.string.hdr."readFile"   �  "go.importpath."".   �  .type.func(*go/ast.File)   �  Ftype.func(*"".reader, *go/ast.File)   �  *"".(*reader).readFile   �  *"".(*reader).readFile   �  0go.string.hdr."readFunc"   �  "go.importpath."".   �  6type.func(*go/ast.FuncDecl)   �  Ntype.func(*"".reader, *go/ast.FuncDecl)   �  *"".(*reader).readFunc   �  *"".(*reader).readFunc   �  0go.string.hdr."readNote"   �  "go.importpath."".   �  8type.func([]*go/ast.Comment)   �  Ptype.func(*"".reader, []*go/ast.Comment)   �  *"".(*reader).readNote   �  *"".(*reader).readNote   �  2go.string.hdr."readNotes"   �  "go.importpath."".   �  Btype.func([]*go/ast.CommentGroup)   �  Ztype.func(*"".reader, []*go/ast.CommentGroup)   �  ,"".(*reader).readNotes   �  ,"".(*reader).readNotes   �  6go.string.hdr."readPackage"   �  "go.importpath."".   �  Ftype.func(*go/ast.Package, "".Mode)   �  ^type.func(*"".reader, *go/ast.Package, "".Mode)   �  0"".(*reader).readPackage   �  0"".(*reader).readPackage   �  0go.string.hdr."readType"   �  "go.importpath."".   �  Xtype.func(*go/ast.GenDecl, *go/ast.TypeSpec)   �  ptype.func(*"".reader, *go/ast.GenDecl, *go/ast.TypeSpec)   �  *"".(*reader).readType   �  *"".(*reader).readType   �  2go.string.hdr."readValue"   �  "go.importpath."".   �  4type.func(*go/ast.GenDecl)   �  Ltype.func(*"".reader, *go/ast.GenDecl)   �  ,"".(*reader).readValue   �  ,"".(*reader).readValue   �  Hgo.string.hdr."recordAnonymousField"   �  "go.importpath."".   �  Xtype.func(*"".namedType, go/ast.Expr) string   �  ptype.func(*"".reader, *"".namedType, go/ast.Expr) string   �  B"".(*reader).recordAnonymousField   �  B"".(*reader).recordAnonymousField   �  0go.string.hdr."remember"   �  "go.importpath."".   �  @type.func(*go/ast.InterfaceType)   �  Xtype.func(*"".reader, *go/ast.InterfaceType)   �  *"".(*reader).remember   �  *"".(*reader).remember   �&runtime.gcbits.cab2   ʲ �4go.string.hdr."doc.reader"             
          ,go.string."doc.reader"   �,go.string."doc.reader"    doc.reader  �(go.string.hdr."mode"                        go.string."mode"   � go.string."mode"   
mode  �2go.string.hdr."filenames"             	          *go.string."filenames"   �*go.string."filenames"    filenames  �*go.string.hdr."notes"                       "go.string."notes"   �"go.string."notes"   notes  �.go.string.hdr."imports"                       &go.string."imports"   �&go.string."imports"   imports  �2go.string.hdr."hasDotImp"             	          *go.string."hasDotImp"   �*go.string."hasDotImp"    hasDotImp  �*go.string.hdr."types"                       "go.string."types"   �"go.string."types"   types  �2go.string.hdr."errorDecl"             	          *go.string."errorDecl"   �*go.string."errorDecl"    errorDecl  �.go.string.hdr."fixlist"                       &go.string."fixlist"   �&go.string."fixlist"   fixlist  �,go.string.hdr."reader"                       $go.string."reader"   �$go.string."reader"   reader  �type."".reader  �  ��       �       ��                                                                                                                                                                                                                     0                                       8                                       @                                       H                                       `                                       h                                       p                                       x                                               T0�  runtime.algarray   @  &runtime.gcbits.cab2   P  4go.string.hdr."doc.reader"   p  type.*"".reader   �� type."".reader   �  (go.string.hdr."mode"   �  "go.importpath."".   �  type."".Mode   �  &go.string.hdr."doc"   �  "go.importpath."".   �  type.string   �  2go.string.hdr."filenames"   �  "go.importpath."".   �  type.[]string   �  *go.string.hdr."notes"   �  "go.importpath."".   �  4type.map[string][]*"".Note   �  .go.string.hdr."imports"   �  "go.importpath."".   �  &type.map[string]int   �  2go.string.hdr."hasDotImp"   �  "go.importpath."".   �  type.bool   �  ,go.string.hdr."values"   �  "go.importpath."".   �   type.[]*"".Value   �  *go.string.hdr."types"   �  "go.importpath."".   �  :type.map[string]*"".namedType   �  *go.string.hdr."funcs"   �  "go.importpath."".   �  "type."".methodSet   �  2go.string.hdr."errorDecl"   �  "go.importpath."".   �  type.bool   �  .go.string.hdr."fixlist"   �  "go.importpath."".   �  8type.[]*go/ast.InterfaceType   `� type."".reader   �  ,go.string.hdr."reader"   �  "go.importpath."".   �� type."".reader   �8go.string.hdr."*doc.Example"                       0go.string."*doc.Example"   �0go.string."*doc.Example"    *doc.Example  � type.*"".Example  �  �              �c4 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  8go.string.hdr."*doc.Example"   p  2go.weak.type.**"".Example   �  type."".Example   �&runtime.gcbits.f504   � �6go.string.hdr."doc.Example"                       .go.string."doc.Example"   �.go.string."doc.Example"    doc.Example  �(go.string.hdr."Code"                        go.string."Code"   � go.string."Code"   
Code  �(go.string.hdr."Play"                        go.string."Play"   � go.string."Play"   
Play  �0go.string.hdr."Comments"                       (go.string."Comments"   �(go.string."Comments"    Comments  �,go.string.hdr."Output"                       $go.string."Output"   �$go.string."Output"   Output  �6go.string.hdr."EmptyOutput"                       .go.string."EmptyOutput"   �.go.string."EmptyOutput"    EmptyOutput  �*go.string.hdr."Order"                       "go.string."Order"   �"go.string."Order"   Order  �type."".Example  �  �p       X       �Hx�                                                                                                                                                                                                                      0                                       8                                       P                                       `                                       h                                               20�  runtime.algarray   @  &runtime.gcbits.f504   P  6go.string.hdr."doc.Example"   p   type.*"".Example   �� type."".Example   �  (go.string.hdr."Name"   �  type.string   �  &go.string.hdr."Doc"   �  type.string   �  (go.string.hdr."Code"   �   type.go/ast.Node   �  (go.string.hdr."Play"   �  "type.*go/ast.File   �  0go.string.hdr."Comments"   �  6type.[]*go/ast.CommentGroup   �  ,go.string.hdr."Output"   �  type.string   �  6go.string.hdr."EmptyOutput"   �  type.bool   �  *go.string.hdr."Order"   �  type.int   `� type."".Example   �  .go.string.hdr."Example"   �  "go.importpath."".   �� type."".Example   �<go.string.hdr."[]*doc.Example"                       4go.string."[]*doc.Example"   �4go.string."[]*doc.Example"    []*doc.Example  �$type.[]*"".Example �  �              B6e[                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."[]*doc.Example"   p  6go.weak.type.*[]*"".Example   �   type.*"".Example   �Pgo.typelink.[]*doc.Example	[]*"".Example              $type.[]*"".Example   �Dgo.string.hdr."*doc.exampleByName"                       <go.string."*doc.exampleByName"   �<go.string."*doc.exampleByName" 0  &*doc.exampleByName  �:go.string.hdr."exampleByName"                       2go.string."exampleByName"   �2go.string."exampleByName"    exampleByName  �&go.string.hdr."Len"                       go.string."Len"   �go.string."Len"   Len  �Tgclocals·33cdeccccebe80329f1fdbee7f5874cb           �Tgclocals·3f5c1f818fa7055d0400cecd34057162             �(go.string.hdr."Swap"                        go.string."Swap"   � go.string."Swap"   
Swap  �Tgclocals·bade3c5f6d433f8d8fecc50019bf4c85                   �Tgclocals·41a13ac73c712c01973b8fe23f62d694                  �(go.string.hdr."Less"                        go.string."Less"   � go.string."Less"   
Less  �Tgclocals·790e5cc5051fc0affc980ade09e929ec              �Tgclocals·2fccd208efe70893f9ac8d682812ae72             �Xgo.string.hdr."func(*doc.exampleByName) int"                       Pgo.string."func(*doc.exampleByName) int"   �Pgo.string."func(*doc.exampleByName) int" @  :func(*doc.exampleByName) int  �@type.func(*"".exampleByName) int �  �              .��A 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."func(*doc.exampleByName) int"   p  Rgo.weak.type.*func(*"".exampleByName) int   �� @type.func(*"".exampleByName) int   �� @type.func(*"".exampleByName) int   �  ,type.*"".exampleByName   �  type.int   ��go.typelink.func(*doc.exampleByName) int	func(*"".exampleByName) int              @type.func(*"".exampleByName) int   �ngo.string.hdr."func(*doc.exampleByName, int, int) bool"             '          fgo.string."func(*doc.exampleByName, int, int) bool"   �fgo.string."func(*doc.exampleByName, int, int) bool" P  Pfunc(*doc.exampleByName, int, int) bool  �Vtype.func(*"".exampleByName, int, int) bool �  �              _H�c 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  ngo.string.hdr."func(*doc.exampleByName, int, int) bool"   p  hgo.weak.type.*func(*"".exampleByName, int, int) bool   �� Vtype.func(*"".exampleByName, int, int) bool   �� Vtype.func(*"".exampleByName, int, int) bool   �  ,type.*"".exampleByName   �  type.int   �  type.int   �  type.bool   ��go.typelink.func(*doc.exampleByName, int, int) bool	func(*"".exampleByName, int, int) bool              Vtype.func(*"".exampleByName, int, int) bool   �dgo.string.hdr."func(*doc.exampleByName, int, int)"             "          \go.string."func(*doc.exampleByName, int, int)"   �\go.string."func(*doc.exampleByName, int, int)" P  Ffunc(*doc.exampleByName, int, int)  �Ltype.func(*"".exampleByName, int, int) �  �              @�g 3                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  dgo.string.hdr."func(*doc.exampleByName, int, int)"   p  ^go.weak.type.*func(*"".exampleByName, int, int)   �� Ltype.func(*"".exampleByName, int, int)   �� Ltype.func(*"".exampleByName, int, int)   �  ,type.*"".exampleByName   �  type.int   �  type.int   ��go.typelink.func(*doc.exampleByName, int, int)	func(*"".exampleByName, int, int)              Ltype.func(*"".exampleByName, int, int)   �4go.string.hdr."func() int"             
          ,go.string."func() int"   �,go.string."func() int"    func() int  �type.func() int �  �              �9� 3                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."func() int"   p  0go.weak.type.*func() int   �� type.func() int   �� type.func() int   �  type.int   �Bgo.typelink.func() int	func() int              type.func() int   �Fgo.string.hdr."func(int, int) bool"                       >go.string."func(int, int) bool"   �>go.string."func(int, int) bool" 0  (func(int, int) bool  �0type.func(int, int) bool �  �              �" 3                                                                                                                    0�  runtime.algarray   @  "runtime.gcbits.01   P  Fgo.string.hdr."func(int, int) bool"   p  Bgo.weak.type.*func(int, int) bool   �� 0type.func(int, int) bool   �� 0type.func(int, int) bool   �  type.int   �  type.int   �  type.bool   �fgo.typelink.func(int, int) bool	func(int, int) bool              0type.func(int, int) bool   �<go.string.hdr."func(int, int)"                       4go.string."func(int, int)"   �4go.string."func(int, int)"    func(int, int)  �&type.func(int, int) �  �              %Ǆ 3                                                                                                              0�  runtime.algarray   @  "runtime.gcbits.01   P  <go.string.hdr."func(int, int)"   p  8go.weak.type.*func(int, int)   �� &type.func(int, int)   �� &type.func(int, int)   �  type.int   �  type.int   �Rgo.typelink.func(int, int)	func(int, int)              &type.func(int, int)   �,type.*"".exampleByName  �  �              �(�� 6                                                                                                                                                                                                                                      ,0�  runtime.algarray   @  "runtime.gcbits.01   P  Dgo.string.hdr."*doc.exampleByName"   p  >go.weak.type.**"".exampleByName   �  *type."".exampleByName   `� ,type.*"".exampleByName   �� ,type.*"".exampleByName   �  &go.string.hdr."Len"   �  type.func() int   �  @type.func(*"".exampleByName) int   �  ."".(*exampleByName).Len   �  ."".(*exampleByName).Len   �  (go.string.hdr."Less"   �  0type.func(int, int) bool   �  Vtype.func(*"".exampleByName, int, int) bool   �  0"".(*exampleByName).Less   �  0"".(*exampleByName).Less   �  (go.string.hdr."Swap"   �  &type.func(int, int)   �  Ltype.func(*"".exampleByName, int, int)   �  0"".(*exampleByName).Swap   �  0"".(*exampleByName).Swap   �Bgo.string.hdr."doc.exampleByName"                       :go.string."doc.exampleByName"   �:go.string."doc.exampleByName" 0  $doc.exampleByName  �Vgo.string.hdr."func(doc.exampleByName) int"                       Ngo.string."func(doc.exampleByName) int"   �Ngo.string."func(doc.exampleByName) int" @  8func(doc.exampleByName) int  �>type.func("".exampleByName) int �  �              %�� 3                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  Vgo.string.hdr."func(doc.exampleByName) int"   p  Pgo.weak.type.*func("".exampleByName) int   �� >type.func("".exampleByName) int   �� >type.func("".exampleByName) int   �  *type."".exampleByName   �  type.int   ��go.typelink.func(doc.exampleByName) int	func("".exampleByName) int              >type.func("".exampleByName) int   �lgo.string.hdr."func(doc.exampleByName, int, int) bool"             &          dgo.string."func(doc.exampleByName, int, int) bool"   �dgo.string."func(doc.exampleByName, int, int) bool" P  Nfunc(doc.exampleByName, int, int) bool  �Ttype.func("".exampleByName, int, int) bool �  �              �iJ� 3                                                                                                                            0�  runtime.algarray   @  "runtime.gcbits.01   P  lgo.string.hdr."func(doc.exampleByName, int, int) bool"   p  fgo.weak.type.*func("".exampleByName, int, int) bool   �� Ttype.func("".exampleByName, int, int) bool   �� Ttype.func("".exampleByName, int, int) bool   �  *type."".exampleByName   �  type.int   �  type.int   �  type.bool   ��go.typelink.func(doc.exampleByName, int, int) bool	func("".exampleByName, int, int) bool              Ttype.func("".exampleByName, int, int) bool   �bgo.string.hdr."func(doc.exampleByName, int, int)"             !          Zgo.string."func(doc.exampleByName, int, int)"   �Zgo.string."func(doc.exampleByName, int, int)" P  Dfunc(doc.exampleByName, int, int)  �Jtype.func("".exampleByName, int, int) �  �              T)�J 3                                                                                                                      0�  runtime.algarray   @  "runtime.gcbits.01   P  bgo.string.hdr."func(doc.exampleByName, int, int)"   p  \go.weak.type.*func("".exampleByName, int, int)   �� Jtype.func("".exampleByName, int, int)   �� Jtype.func("".exampleByName, int, int)   �  *type."".exampleByName   �  type.int   �  type.int   ��go.typelink.func(doc.exampleByName, int, int)	func("".exampleByName, int, int)              Jtype.func("".exampleByName, int, int)   �*type."".exampleByName  �  �              3��                                                                                                                                                                                                                                       00�  runtime.algarray   @  "runtime.gcbits.01   P  Bgo.string.hdr."doc.exampleByName"   p  ,type.*"".exampleByName   �   type.*"".Example   `� *type."".exampleByName   �  :go.string.hdr."exampleByName"   �  "go.importpath."".   �� *type."".exampleByName   �  &go.string.hdr."Len"   �  type.func() int   �  >type.func("".exampleByName) int   �  ."".(*exampleByName).Len   �  ("".exampleByName.Len   �  (go.string.hdr."Less"   �  0type.func(int, int) bool   �  Ttype.func("".exampleByName, int, int) bool   �  0"".(*exampleByName).Less   �  *"".exampleByName.Less   �  (go.string.hdr."Swap"   �  &type.func(int, int)   �  Jtype.func("".exampleByName, int, int)   �  0"".(*exampleByName).Swap   �  *"".exampleByName.Swap   �6go.string.hdr."[]*ast.File"                       .go.string."[]*ast.File"   �.go.string."[]*ast.File"    []*ast.File  �&type.[]*go/ast.File �  �              ��=s                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  6go.string.hdr."[]*ast.File"   p  8go.weak.type.*[]*go/ast.File   �  "type.*go/ast.File   �Lgo.typelink.[]*ast.File	[]*go/ast.File              &type.[]*go/ast.File   �4go.string.hdr."[]ast.Decl"             
          ,go.string."[]ast.Decl"   �,go.string."[]ast.Decl"    []ast.Decl  �$type.[]go/ast.Decl �  �              q|�+                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."[]ast.Decl"   p  6go.weak.type.*[]go/ast.Decl   �   type.go/ast.Decl   �Hgo.typelink.[]ast.Decl	[]go/ast.Decl              $type.[]go/ast.Decl   �4go.string.hdr."**ast.File"             
          ,go.string."**ast.File"   �,go.string."**ast.File"    **ast.File  �$type.**go/ast.File �  �              Q�I� 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  4go.string.hdr."**ast.File"   p  6go.weak.type.***go/ast.File   �  "type.*go/ast.File   �:go.string.hdr."[]*ast.Object"                       2go.string."[]*ast.Object"   �2go.string."[]*ast.Object"    []*ast.Object  �*type.[]*go/ast.Object �  �              �.H�                                                 
0�  runtime.algarray   @  "runtime.gcbits.01   P  :go.string.hdr."[]*ast.Object"   p  <go.weak.type.*[]*go/ast.Object   �  &type.*go/ast.Object   �Tgo.typelink.[]*ast.Object	[]*go/ast.Object              *type.[]*go/ast.Object   �<go.string.hdr."[8]*ast.Object"                       4go.string."[8]*ast.Object"   �4go.string."[8]*ast.Object"    [8]*ast.Object  �,type.[8]*go/ast.Object �  �@       @       7˂4                                                                0  type..alg64   @  "runtime.gcbits.ff   P  <go.string.hdr."[8]*ast.Object"   p  >go.weak.type.*[8]*go/ast.Object   �  &type.*go/ast.Object   �  *type.[]*go/ast.Object   �Xgo.typelink.[8]*ast.Object	[8]*go/ast.Object              ,type.[8]*go/ast.Object   �Xgo.string.hdr."*map.bucket[*ast.Object]bool"                       Pgo.string."*map.bucket[*ast.Object]bool"   �Pgo.string."*map.bucket[*ast.Object]bool" @  :*map.bucket[*ast.Object]bool  �Htype.*map.bucket[*go/ast.Object]bool �  �              V�_l 6                                                
0�  runtime.algarray   @  "runtime.gcbits.01   P  Xgo.string.hdr."*map.bucket[*ast.Object]bool"   p  Zgo.weak.type.**map.bucket[*go/ast.Object]bool   �  Ftype.map.bucket[*go/ast.Object]bool   �Vgo.string.hdr."map.bucket[*ast.Object]bool"                       Ngo.string."map.bucket[*ast.Object]bool"   �Ngo.string."map.bucket[*ast.Object]bool" @  8map.bucket[*ast.Object]bool  �Ftype.map.bucket[*go/ast.Object]bool �  �X       X       `Q�C                                                                                                                                                                              H                                       P       0�  runtime.algarray   @  &runtime.gcbits.fe05   P  Vgo.string.hdr."map.bucket[*ast.Object]bool"   p  Xgo.weak.type.*map.bucket[*go/ast.Object]bool   �� Ftype.map.bucket[*go/ast.Object]bool   �  .go.string.hdr."topbits"   �  type.[8]uint8   �  (go.string.hdr."keys"   �  ,type.[8]*go/ast.Object   �  ,go.string.hdr."values"   �  type.[8]bool   �  0go.string.hdr."overflow"   �  Htype.*map.bucket[*go/ast.Object]bool   �Pgo.string.hdr."map.hdr[*ast.Object]bool"                       Hgo.string."map.hdr[*ast.Object]bool"   �Hgo.string."map.hdr[*ast.Object]bool" @  2map.hdr[*ast.Object]bool  �@type.map.hdr[*go/ast.Object]bool � 